H   ����@        ����@����@����@                ����@����@H                     x   �\�qMY�p�O�A�-�.�����L�r������p���Im�O�:�}j��$�7�оg�ƾ7�о�$�}j�O�:��Im��p�����r�࿊L����-�.�A�p�O�qMY�x   x   qMY�g�R�W�F�k6��:#�&�� ��xʿ����!��e�P�$�q�#�۾�Ǿ�Ǿ&�۾r�$�^�P��!������xʿ��&���:#�~k6�V�F�h�R�pMY�x   x   p�O�W�F��9���'�mb�' �,�׿N��2ُ��d���3��R�m`��Wʾ�����Wʾq`辂R���3�y�d�/ُ�M��,�׿' �nb���'��9�W�F�r�O�h�R�x   x   A�k6���'�	g���L��R�� �ou�a�A�!���$��`�ξ�绾�绾f�ξ�$��#��\�A�nu� �R��Q��	��g���'�k6�A�W�F�V�F�x   x   -�.��:#�mb����{㿫$�������q��ڍL���!��u �F`Ӿ�&��R����&��@`Ӿ�u ���!��L��q�������$���{���pb��:#�-�.�k6��9�~k6�x   x   ���&��' �L�࿫$��\���H����jS� �'�P5�(�׾Bط�`5��f5��@ط�2�׾R5�%�'��jS�F���\����$��O��( �%������:#���'���'��:#�x   x   �L� ��,�׿R������H���{�U�E++�J���۾�o���l��Rz���l���o����۾J�E++�~�U�I�������R��-�׿��L�%��pb�g�nb�&��x   x   r�࿷xʿN�� 𘿬q���jS�E++�k[	���ݾ~l���מ�J���O����מ�|l����ݾh[	�H++��jS��q��!�K���xʿr����( ���	��' ���x   x   ������2ُ�ou�ڍL� �'�J���ݾ'v���$��߭��Q���ݭ���$��(v����ݾJ�%�'��L�ju�/ُ��������xʿ-�׿O�࿛{�Q��,�׿�xʿx   x   �p���!���d�a�A���!�P5���۾~l���$�����9���8�������$��l����۾O5���!�`�A���d��!���p�����K��R���$���$��R��M�����x   x   �Im�e�P���3�!���u �(�׾�o���מ�߭��9���vG��>���᭍��מ��o��(�׾�u �#����3�_�P��Im��!��/ُ�!�����\������� �/ُ��!��x   x   O�:�$��R��$��F`ӾBط��l��J���Q���8���>���L���M����l��6ط�X`Ӿ�$���R�$�G�:�_�P���d�ju��q��I���F����q��nu�y�d�^�P�x   x   }j�q�m`�`�ξ�&��`5��Rz��O���ݭ�����᭍�M���Kz��[5���&��o�ξn`�p�tj�$���3�`�A��L��jS�~�U��jS��L�\�A���3�$�x   x   �$�#�۾�Wʾ�绾R���f5���l���מ��$���$���מ��l��[5��a����绾�Wʾ%�۾�$�p��R�#����!�%�'�H++�E++�%�'���!�#���R�r�x   x   7�о�Ǿ�����绾�&��@ط��o��|l��(v��l���o��6ط��&���绾�����Ǿ1�о%�۾n`辣$���u �O5�J�h[	�J�R5��u ��$��q`�&�۾x   x   g�ƾ�Ǿ�Wʾf�ξ@`Ӿ2�׾��۾��ݾ��ݾ��۾(�׾X`Ӿo�ξ�Wʾ�Ǿ\�ƾ�Ǿ�Wʾo�ξX`Ӿ(�׾��۾��ݾ��ݾ��۾2�׾@`Ӿf�ξ�Wʾ�Ǿx   x   7�о&�۾q`辠$���u �R5�J�h[	�J�O5��u ��$��n`�%�۾1�о�Ǿ�����绾�&��6ط��o��l��(v��|l���o��@ط��&���绾�����Ǿx   x   �$�r��R�#����!�%�'�E++�H++�%�'���!�#���R�p��$�%�۾�Wʾ�绾a���[5���l���מ��$���$���מ��l��f5��R����绾�Wʾ#�۾x   x   }j�$���3�\�A��L��jS�~�U��jS��L�`�A���3�$�tj�p�n`�o�ξ�&��[5��Kz��M���᭍����ݭ��O���Rz��`5���&��`�ξm`�q�x   x   O�:�^�P�y�d�nu��q��F���I����q��ju���d�_�P�G�:�$��R��$��X`Ӿ6ط��l��M���L���>���8���Q���J����l��Bط�F`Ӿ�$���R�$�x   x   �Im��!��/ُ� �����\�������!�/ُ��!���Im�_�P���3�#���u �(�׾�o���מ�᭍�>���vG��9���߭���מ��o��(�׾�u �!����3�e�P�x   x   �p�����M��R���$���$��R��K������p���!����d�`�A���!�O5���۾l���$�����8���9�������$��~l����۾P5���!�a�A��d��!��x   x   ����xʿ,�׿Q�࿛{�O��-�׿�xʿ������/ُ�ju��L�%�'�J���ݾ(v���$��ݭ��Q���߭���$��'v����ݾJ� �'�ڍL�ou�2ُ����x   x   r����' �	����( ���r�࿹xʿK��!𘿭q���jS�H++�h[	���ݾ|l���מ�O���J����מ�~l����ݾk[	�E++��jS��q�� �N���xʿx   x   �L�&��nb�g�pb�%���L���-�׿R������I���~�U�E++�J���۾�o���l��Rz���l���o����۾J�E++�{�U�H�������R��,�׿ ��x   x   ����:#���'���'��:#����%��( �O�࿨$��\���F����jS�%�'�R5�2�׾@ط�f5��`5��Bط�(�׾P5� �'��jS�H���\����$��L��' �&��x   x   -�.�~k6��9�k6�-�.��:#�pb����{㿪$�������q���L���!��u �@`Ӿ�&��R����&��F`Ӿ�u ���!�ڍL��q�������$���{���mb��:#�x   x   A�V�F�W�F�A�k6���'�g�	��Q��R�� �nu�\�A�#���$��f�ξ�绾�绾`�ξ�$��!��a�A�ou� �R��L����	g���'�k6�x   x   p�O�h�R�r�O�W�F��9���'�nb�' �,�׿M��/ُ�y�d���3��R�q`��Wʾ�����Wʾm`辀R���3��d�2ُ�N��,�׿' �mb���'��9�W�F�x   x   qMY�pMY�h�R�V�F�~k6��:#�&����xʿ����!��^�P�$�r�&�۾�Ǿ�Ǿ#�۾q�$�e�P��!������xʿ ��&���:#�k6�W�F�g�R�x   x   qMY�g�R�W�F�k6��:#�&�� ��xʿ����!��e�P�$�q�#�۾�Ǿ�Ǿ&�۾r�$�^�P��!������xʿ��&���:#�~k6�V�F�h�R�pMY�x   x   g�R��I�m�;� *�&g�|����ڿd\��٪��=cg�6������-V̾={¾(V̾������6�Hcg�ߪ��f\����ڿz��&g�*�m�;��I�h�R���U�x   x   W�F�m�;�},�̈�j�6}�2���؜�\7{�xF��Q�w���Ҿs��s���Ҿw���Q�xF�\7{��؜�2��2}�j�͈�},�n�;�U�F���L���L�x   x   k6� *�̈������`�ǿ�Ӥ��L��oT��;'�H����پ3I��uX��1I����پF���;'�tT��L���Ӥ�`�ǿ�����͈� *�k6�ZX>�aA�[X>�x   x   �:#�&g�j����Eʿt���(-����]�3�/���B��}r��gޭ�iޭ�yr��H�ྏ�1�/���]�$-��v����Eʿ��k�&g��:#��,��_1��_1��,�x   x   &��|��6}�`�ǿt����؋���b�l95�
���c�BR��&����<��$���?R���c���h95���b��؋�t���e�ǿ5}�x��'��uw�o��!�o��sw�x   x    ���ڿ2���Ӥ�(-����b�N7�9��<꾈O��hj��<:��=:��lj���O���<�9�M7���b�'-���Ӥ�2����ڿ����p�
�ǂ�Ȃ�r�
���x   x   �xʿd\���؜��L����]�l95�9����q���ʠ��*w��eΌ�,w��Ϡ��u������9�g95���]��L���؜�d\���xʿ~�ݿ���2���u���2����}�ݿx   x   ���٪��\7{�oT�3�/�
���<�q���Q��⩏�[��\��穏�V��v����<���0�/�lT�W7{�ݪ�����i����Mſ@�Ͽ�$տ�$տ@�Ͽ�Mſk���x   x   �!��=cg�xF��;'����c澈O��ʠ��⩏�/郾���0郾婏�Ǡ���O���c澑��;'�xF�Ccg��!����������^��P���g8��O����^���������x   x   e�P�6��Q�H��B��BR��hj��*w��[��������W��1w��jj��GR��F��A���Q�6�g�P��_j�d���ň���m�������m��È��f����_j�x   x   $���w����پ}r��&���<:��eΌ�\��0郾W��fΌ�@:��0����r����پw�����$��]8���K�L\��Ki��q�d]t��q��Ki�L\���K��]8�x   x   q�����Ҿ3I��gޭ��<��=:��,w��穏�婏�1w��@:���<��jޭ�I���Ҿ���u�!���> ���-���8�ީ@���D���D�ک@���8���-��> ���x   x   #�۾-V̾s��uX��iޭ�$���lj��Ϡ��V��Ǡ��jj��0���jޭ�fX��s��3V̾%�۾���W? ��	���f��l��n4�l��d������	�V? ����x   x   �Ǿ={¾s��1I��yr��?R���O��u���v����O��GR���r��I��s��C{¾�Ǿ`�ξq׾;5���꾒�����Bb��Vb������������<5�q׾Y�ξx   x   �Ǿ(V̾�Ҿ��پH���c��<�����<��c�F�ྗ�پ�Ҿ3V̾�ǾȠľ��þ2�ľ�ƾ�`ɾ�˾�;x�ξ#�;��˾�`ɾ$�ƾ3�ľ��þ��ľx   x   &�۾���w��F������9�9�����A��w�����%�۾`�ξ��þU4��"���������R���Ȭ��Ȭ�R���������,��N4����þY�ξx   x   r�����Q��;'�1�/�h95�M7�g95�0�/��;'��Q����u����q׾2�ľ"��b
��e@��p[��R�������Y���f[��T@��f
��5��4�ľq׾���x   x   $�6�xF�tT���]���b���b���]�lT�xF�6�$�!��W? �;5��ƾ���e@�����[7���^���^��_7�����Z@�����%�ƾ35�Z? ���x   x   ^�P�Hcg�\7{��L��$-���؋�'-���L��W7{�Ccg�g�P��]8��> ��	���꾼`ɾ����p[��[7����5���Z7��e[�������`ɾ�����	��> ��]8�x   x   �!��ߪ���؜��Ӥ�v���t����Ӥ��؜�ݪ���!���_j���K���-�������˾R��R����^���5���5���^��Y���R����˾�������-���K��_j�x   x   ���f\��2��`�ǿ�Eʿe�ǿ2��d\��������d���L\���8�f�������;�Ȭ������^����^�������Ȭ��;����l����8�L\�a������x   x   �xʿ��ڿ2}�����5}濑�ڿ�xʿi�������ň���Ki�ީ@�l��Bb��x�ξ�Ȭ�Y���_7��Z7��Y����Ȭ�v�ξHb��l���@��Ki�ƈ������k���x   x   ��z��j����k�x����~�ݿ�Mſ�^���m���q���D�n4�Vb��#�;R��f[�����e[��R���;Hb��v4���D��q��m���^���Mſ}�ݿx   x   &��&g�͈�͈�&g�'������@�ϿP�����d]t���D�l��������˾����T@��Z@��������˾����l����D�^]t���N���@�Ͽ����x   x   �:#�*�},� *��:#�uw�p�
��2���$տg8�����q�ک@�d������`ɾ���f
������`ɾ���l���@��q���e8���$տ�2��s�
�sw�x   x   ~k6�m�;�n�;�k6��,�o��ǂ��u���$տO����m���Ki���8������$�ƾ,��5��%�ƾ�������8��Ki��m��N����$տ�u��Ȃ�n���,�x   x   V�F��I�U�F�ZX>��_1�!�Ȃ��2��@�Ͽ�^��È��L\���-���	�<5�3�ľN4��4�ľ35���	���-�L\�ƈ���^��@�Ͽ�2��Ȃ�!��_1�[X>�x   x   h�R�h�R���L�aA��_1�o��r�
��쿟Mſ����f�����K��> �V? �q׾��þ��þq׾Z? ��> ���K�a��������Mſ��s�
�n���_1�`A���L�x   x   pMY���U���L�[X>��,�sw���}�ݿk�������_j��]8������Y�ξ��ľY�ξ������]8��_j����k���}�ݿ��sw��,�[X>���L���U�x   x   p�O�W�F��9���'�mb�' �,�׿N��2ُ��d���3��R�m`��Wʾ�����Wʾq`辂R���3�y�d�/ُ�M��,�׿' �nb���'��9�W�F�r�O�h�R�x   x   W�F�m�;�},�̈�j�6}�2���؜�\7{�xF��Q�w���Ҿs��s���Ҿw���Q�xF�\7{��؜�2��2}�j�͈�},�n�;�U�F���L���L�x   x   �9�},���c�
���;JʿY�����0�V�00)�_+�2�۾�
�������
��;�۾b+�10)�!�V�����Y�=Jʿ��b�
���},��9�aA�_�C�`A�x   x   ��'�̈�c�
�m�� �ϿnP�������:c�:�3�J.�C�H����а��а�I���?�L.�9�3��:c�����lP��!�Ͽl��c�
�͈���'��_1�rl6�pl6��_1�x   x   mb�j��� �Ͽ������L3k�j�;����C�-Wľ̮���椾̮��3Wľ�C���h�;�H3k�������"�Ͽ��i�ob�n���~%���'��~%�n��x   x   ' �6}�;JʿnP������m�L�?�t��Z��ƾ&��,��,��&���ƾ&Z�z��S�?���m���lP��;Jʿ6}�( �r�
� h�bj�`j�h�s�
�x   x   ,�׿2��Y�����L3k�L�?�_��י��LjȾ�è�`J��q-��[J���è�QjȾݙ��Z��M�?�B3k�����W�2��1�׿�쿯���و�;K�׈�������x   x   N���؜������:c�j�;�t��י���ɾ,��K钾�j���j��I钾
,���ɾԙ��v��o�;��:c������؜�N���Mſ�6տؗ�����՗��6տ�Mſx   x   2ُ�\7{�0�V�:�3���Z�LjȾ,��Fϑ�����mG������?ϑ�	,��MjȾZ���;�3�)�V�[7{�1ُ�����xׯ�ba���¿�3ſ�¿ea��vׯ�����x   x   �d�xF�00)�J.��C��ƾ�è�K钾����P1{�J1{�����H钾�è��ƾ�C�N.�/0)�xF�w�d�b���������cˠ��٤��٤�cˠ�������a���x   x   ��3��Q�_+�C�-Wľ&��`J���j��mG��J1{�qG���j��WJ��&��&WľE�d+��Q���3���K� �a��;u��!���䆿!����䆿�!���;u� �a���K�x   x   �R�w��2�۾H���̮��,��q-���j�����������j��j-��,��Ǯ��J���J�۾w���R��> ���1���A��9O�d�X��]��]�b�X��9O���A���1��> �x   x   m`��Ҿ�
���а��椾,��[J��I钾?ϑ�H钾WJ��,���椾�а��
���Ҿf`�U? ���������#���+� M1�x!3��L1���+���#�������Z? �x   x   �Wʾs�������а�̮��&���è�
,��	,���è�&��Ǯ���а�����s���Wʾ	q׾�#�y��v�PU�����N��N����OU�u�y���#�q׾x   x   ����s���
��I���3Wľ�ƾQjȾ�ɾMjȾ�ƾ&WľJ����
��s��������þȾ��ξF�վܾ߯�_⾤&�Oy羝&澒_��ܾB�վ��ξɏȾ��þx   x   �Wʾ�Ҿ;�۾?徢C�&Z�ݙ��ԙ��Z�C�E�J�۾�Ҿ�Wʾ��þ=���=���D��茻�~��у��'��'��΃��~��ڌ���D��=��A�����þx   x   q`�w��b+�L.���z��Z��v����N.�d+�w��f`�	q׾Ⱦ=������&t��e���Hj��(����0��.���[j��]���t������=��ɏȾq׾x   x   �R��Q�10)�9�3�h�;�S�?�M�?�o�;�;�3�/0)��Q��R�U? ��#澐�ξ�D��&t���G��h������\���\����o����G��t���D����ξ�#�V? �x   x   ��3�xF�!�V��:c�H3k���m�B3k��:c�)�V�xF���3��> ����y��F�վ茻�e���h���N�������������Q���t���^���،��B�վ�x������> �x   x   y�d�\7{���������������������[7{�w�d���K���1����v�ܾ߯~��Hj��������v~��v~������Vj��~��دܾw������1���K�x   x   /ُ��؜�Y�lP������lP��W��؜�1ُ�b��� �a���A���#�PU��_�у��(����\�������v~������\��3���ك���_�LU���#���A� �a�f���x   x   M��2��=Jʿ!�Ͽ"�Ͽ;Jʿ2��N����������;u��9O���+�����&�'���0���\���������\���0��'���&澬����+��9O��;u��������x   x   ,�׿2}���l����6}�1�׿�Mſxׯ�����!��d�X� M1��N�Oy�'��.�����Q�����3���'��Ly��N��L1�`�X��!�����vׯ��Mſx   x   ' �j�b�
�c�
�i�( ����6տba��cˠ��䆿�]�x!3��N��&�΃��[j��o���t���Vj��ك���&��N�x!3��]��䆿aˠ�ga���6տ��x   x   nb�͈���͈�ob�r�
�����ؗ��¿�٤�!����]��L1�����_�~��]����G��^���~���_⾬���L1��]�����٤��¿ח࿲���r�
�x   x   ��'�},�},���'�n�� h�و��濂3ſ�٤��䆿b�X���+�OU��ܾڌ��t��t��،��دܾLU���+�`�X��䆿�٤��3ſ��ֈ�h�o��x   x   �9�n�;��9��_1��~%�bj�;K����¿cˠ��!���9O���#�u�B�վ�D�������D��B�վw���#��9O��!��aˠ��¿��;K�`j��~%��_1�x   x   W�F�U�F�aA�rl6���'�`j�׈�՗�ea������;u���A����y����ξ=��=����ξ�x�������A��;u����ga��ח�ֈ�`j���'�pl6�aA�x   x   r�O���L�_�C�pl6��~%�h������6տvׯ���� �a���1�����#�ɏȾA���ɏȾ�#������1� �a����vׯ��6տ����h��~%�pl6�_�C���L�x   x   h�R���L�`A��_1�n��s�
��쿜Mſ����a�����K��> �Z? �q׾��þ��þq׾V? ��> ���K�f��������Mſ��r�
�o���_1�aA���L�h�R�x   x   A�k6���'�	g���L��R�� �ou�a�A�!���$��`�ξ�绾�绾f�ξ�$��#��\�A�nu� �R��Q��	��g���'�k6�A�W�F�V�F�x   x   k6� *�̈������`�ǿ�Ӥ��L��oT��;'�H����پ3I��uX��1I����پF���;'�tT��L���Ӥ�`�ǿ�����͈� *�k6�ZX>�aA�[X>�x   x   ��'�̈�c�
�m�� �ϿnP�������:c�:�3�J.�C�H����а��а�I���?�L.�9�3��:c�����lP��!�Ͽl��c�
�͈���'��_1�rl6�pl6��_1�x   x   	g����m���=ҿ仱�쒿gn��=��$����Cƾ����(�����>ƾ{���$�#�=�rn�쒿仱��=ҿm�����	g�!���'�� *���'�!�x   x   ���� �Ͽ仱�3���ɭs�+D�V��w ��ʾ�����=���=������ʾr ��Q��(D���s�6���滱�!�Ͽ����Ȃ�aj�Ս�Ս�`j�Ȃ�x   x   L��`�ǿnP��쒿ɭs��2F����1���
7;b����[���Z��7;,�������2F�ʭs�쒿nP��a�ǿN���2��ֈ����H�
����ֈ��2��x   x   R���Ӥ�����gn�+D���������ξT﫾wS��0-��2-��yS��N﫾��ξ������(D�on������Ӥ�R��>�Ͽۗ࿏�쿨���򿍫�ח�@�Ͽx   x    ��L���:c��=�V��1�����ξ$�U����f�� ����f��U���'���ξ=���U���=��:c��L��!��^��ga��v�ǿ��Ͽcҿ��Ͽv�ǿga���^��x   x   ou�oT�:�3��$�w ��
7;T﫾U���5Ճ��x��x�4Ճ�^���N﫾7;l ���$�:�3�wT�pu�È�������nz��<뱿=뱿nz���󤿫��ƈ��x   x   a�A��;'�J.����ʾb��wS���f���x� �q��x��f��zS��^��ʾx��I.��;'�^�A�L\��;u��p��ԍ�@$��,���C$��ԍ��p���;u�L\�x   x   !��H��C�Cƾ�����0-�� ����x��x�����2-�������Hƾ<�H��"����-���A��`T�b�c�׉n�7t�7t�։n�]�c��`T���A���-�x   x   �$����پH�������=���[��2-���f��4Ճ��f��2-���[���=�����C�����پ�$����	������'��X4�P>���D�y�F���D�P>��X4���'������	�x   x   `�ξ3I���а��(���=���yS��U���^���zS����=���(���а�I��k�ξ@5��x��7���C����2��4����>�� ��2��x��35�x   x   �绾uX���а��������Z��N﫾'�N﫾^����������а�hX���绾8�ľ��ξ�^ھ��+��gw�����څ ����hw��&���}^ھ��ξ4�ľx   x   �绾1I��I���>ƾʾ7;��ξ��ξ7;ʾHƾC���I���绾T4��	=���ﾾ��¾�@Ǿ�s˾��ξ�о�о��ξ�s˾�@Ǿ��¾�ﾾ=��N4��x   x   f�ξ��پ?�{��r ��,������=���l ��x��<從�پk�ξ8�ľ	=�������±�`@�����'�������옭�����-������a@��ñ�����=��3�ľx   x   �$��F��L.��$�Q��������U���$�I.�H���$��@5ᾊ�ξ�ﾾ�±��\�������V������l���l�����V�������\���±��ﾾ��ξ<5�x   x   #���;'�9�3�#�=�(D��2F�(D��=�:�3��;'�"����	��x���^ھ��¾`@��������G㋾�.������.��B㋾�򓾴���`@����¾}^ھy����	�x   x   \�A�tT��:c�rn���s�ʭs�on��:c�wT�^�A���-����7����@Ǿ����V��G㋾΀��!�{��{�ـ��B㋾�V������@Ǿ�2������-�x   x   nu��L������쒿6���쒿�����L��pu�L\���A���'���+��s˾'�������.��!�{���u��{��.��{��,����s˾1�� ����'���A�L\�x   x    ��Ӥ�lP��仱�滱�nP���Ӥ�!�È���;u��`T��X4�C��gw����ξ�����l������{��{�%����l��������ξlw��B���X4��`T��;u�È��x   x   R��`�ǿ!�Ͽ�=ҿ!�Ͽa�ǿR���^������p��b�c�P>�������о옭��l���.��ـ���.���l��瘭��о�����P>�f�c��p������^��x   x   Q����l��m����N��>�Ͽga����ԍ�׉n���D�2��څ ��о������B㋾B㋾{�������оޅ �4����D�։n�ԍ���ea��@�Ͽx   x   	�����c�
�������2��ۗ�v�ǿnz��@$��7t�y�F�4�������ξ-����V�����V��,�����ξ���4��z�F�7t�C$��oz��v�ǿ՗��2��x   x   g�͈�͈�	g�Ȃ�ֈ���쿳�Ͽ<뱿,���7t���D���hw���s˾���������������s˾lw������D�7t�)���=뱿��Ͽ���׈�Ȃ�x   x   ��'� *���'�!�aj�������cҿ=뱿C$��׉n�P>�>��&���@Ǿa@���\��`@���@Ǿ1��B��P>�։n�C$��=뱿cҿ�����`j�!�x   x   k6�k6��_1���'�Ս�H�
���򿶯Ͽnz��ԍ�]�c��X4� ��澓�¾ñ��±���¾� ���X4�f�c�ԍ�oz����Ͽ���J�
�Ս���'��_1�x   x   A�ZX>�rl6�� *�Ս�������v�ǿ�󤿍p���`T���'�2�}^ھ�ﾾ�����ﾾ}^ھ2���'��`T��p����v�ǿ��쿪��Ս�� *�rl6�ZX>�x   x   W�F�aA�pl6���'�`j�ֈ�ח�ga������;u���A�����x����ξ=��=����ξy�������A��;u����ea��՗�׈�`j���'�rl6�aA�U�F�x   x   V�F�[X>��_1�!�Ȃ��2��@�Ͽ�^��ƈ��L\���-���	�35�4�ľN4��3�ľ<5���	���-�L\�È���^��@�Ͽ�2��Ȃ�!��_1�ZX>�U�F��I�x   x   -�.��:#�mb����{㿫$�������q��ڍL���!��u �F`Ӿ�&��R����&��@`Ӿ�u ���!��L��q�������$���{���pb��:#�-�.�k6��9�~k6�x   x   �:#�&g�j����Eʿt���(-����]�3�/���B��}r��gޭ�iޭ�yr��H�ྏ�1�/���]�$-��v����Eʿ��k�&g��:#��,��_1��_1��,�x   x   mb�j��� �Ͽ������L3k�j�;����C�-Wľ̮���椾̮��3Wľ�C���h�;�H3k�������"�Ͽ��i�ob�n���~%���'��~%�n��x   x   ���� �Ͽ仱�3���ɭs�+D�V��w ��ʾ�����=���=������ʾr ��Q��(D���s�6���滱�!�Ͽ����Ȃ�aj�Ս�Ս�`j�Ȃ�x   x   �{��Eʿ����3���7�v��tH��� ��	 ���ξ5����������5����ξ�	 ��� ��tH�F�v�1��������Eʿ�{��u��<K�I�
�A��J�
�;K��u��x   x   �$��t�����ɭs��tH�x6"��"��ҾO����.!��/!������S�Ҿ�"�w6"��tH���s���u����$���$տ�濧��!w��!w��������$տx   x   ����(-��L3k�+D��� ��"�7.Ӿg������� ������ ������ g��;.Ӿ�"��� �*D�P3k�'-�� ���M����¿��ϿF�׿O�ڿH�׿��Ͽ�¿N���x   x   �q����]�j�;�V���	 ��Ҿg���s������W[v�V[v������s��g���Ҿ|	 �U��h�;���]��q���m��cˠ�nz��N����?���?��M���oz��aˠ��m��x   x   ڍL�3�/���w ����ξO��������Pwr���k�Uwr���������P��ξ} ����0�/�ݍL��Ki��!��ԍ��䖿���b�������䖿ԍ��!���Ki�x   x   ��!����C�ʾ5������� ��W[v���k���k�T[v�� ������5��ʾ�C��}�!���8��9O�g�c��~t�_B���c���c��`B���~t�f�c��9O���8�x   x   �u �B��-Wľ�������.!�����V[v�Uwr�T[v����.!���������+WľI���u �����#��X4���B��BN�YqU��W�VqU��BN���B��X4���#���x   x   F`Ӿ}r��̮���=����/!��� ����������� ��.!�����=��®���r��Q`Ӿ���x�!���5�=�#���*��c.��c.���*�=�#��5� ��w����x   x   �&��gޭ��椾�=��������������s��������������=���椾qޭ��&���ƾA�վ��0���(�R���x�����x�Q��(�=����B�վ%�ƾx   x   R���iޭ�̮������5��S g��g��P5������®��qޭ�`���'���D����¾%˾�\ӾA�ھ�߾�������߾:�ھ�\Ӿ%˾��¾�D��5��x   x   �&��yr��3Wľʾ��ξ�Ҿ;.Ӿ�Ҿ��ξʾ+Wľ�r���&��'�������±��j������P��2k��빾�u��빾$k���P������j���±�����,��x   x   @`ӾH�ྡྷC�r ���	 ��"��"�|	 �} ���C�I��Q`Ӿ�ƾ�D���±��M��	褾�?���������-��-��
��������?���社�M��ñ��D��$�ƾx   x   �u �����Q���� �w6"��� �U�������u ����A�վ��¾�j��	褾�H���x���+�����������+���x���H��	褾�j����¾B�վ���x   x   ��!�1�/�h�;�(D��tH��tH�*D�h�;�0�/�}�!���x���%˾����?���x�������E�z�A�z�����𷇾�x���?�����%˾�u���x   x   �L���]�H3k���s�F�v���s�P3k���]�ݍL���8���#�!��0����\Ӿ�P�������+��������r���m���r������+�������P���\Ӿ=��� ����#���8�x   x   �q��$-����6���1�����'-���q���Ki��9O��X4��5�(�A�ھ2k��������E�z���m���m�=�z�������'k��D�ھ(��5��X4��9O��Ki�x   x   ����v�������滱�����u��� ����m���!��g�c���B�=�#�R���߾빾-����A�z���r�=�z���-��#빾�߾T��:�#���B�]�c��!���m��x   x   �$���Eʿ"�Ͽ!�Ͽ�Eʿ�$��M���cˠ�ԍ��~t��BN���*��x�����u��-����������������-���u�����~x���*��BN��~t�ԍ�bˠ�O���x   x   �{������쿜{��$տ�¿nz���䖿_B��YqU��c.�������빾
����+��𷇾�+�����#빾��⾮���c.�YqU�^B���䖿nz���¿�$տx   x   ��k�i����u���濰�ϿN�������c���W��c.��x��߾$k�������x���x������'k���߾~x��c.�t�W��c�����M�����Ͽ���u��x   x   pb�&g�ob�Ȃ�<K����F�׿�?��b����c��VqU���*�Q��:�ھ�P���?���H���?���P��D�ھT����*�YqU��c��_����?��H�׿���;K�ǂ�x   x   �:#��:#�n��aj�I�
�!w��O�ڿ�?�����`B���BN�=�#�(��\Ӿ����社	褾����\Ӿ(�:�#��BN�^B������?��R�ڿ!w��H�
�bj�o��x   x   -�.��,��~%�Ս�A��!w��H�׿M����䖿�~t���B��5�=���%˾�j���M���j��%˾=����5���B��~t��䖿M���H�׿!w��A��Ս��~%��,�x   x   k6��_1���'�Ս�J�
���򿯯Ͽoz��ԍ�f�c��X4� ��澖�¾�±�ñ���¾� ���X4�]�c�ԍ�nz����Ͽ���H�
�Ս���'��_1�k6�x   x   �9��_1��~%�`j�;K����¿aˠ��!���9O���#�w�B�վ�D�������D��B�վu���#��9O��!��bˠ��¿��;K�bj��~%��_1��9�n�;�x   x   ~k6��,�n��Ȃ��u���$տN����m���Ki���8������%�ƾ5��,��$�ƾ�������8��Ki��m��O����$տ�u��ǂ�o���,�k6�n�;�m�;�x   x   ���&��' �L�࿫$��\���H����jS� �'�P5�(�׾Bط�`5��f5��@ط�2�׾R5�%�'��jS�F���\����$��O��( �%������:#���'���'��:#�x   x   &��|��6}�`�ǿt����؋���b�l95�
���c�BR��&����<��$���?R���c���h95���b��؋�t���e�ǿ5}�x��'��uw�o��!�o��sw�x   x   ' �6}�;JʿnP������m�L�?�t��Z��ƾ&��,��,��&���ƾ&Z�z��S�?���m���lP��;Jʿ6}�( �r�
� h�bj�`j�h�s�
�x   x   L��`�ǿnP��쒿ɭs��2F����1���
7;b����[���Z��7;,�������2F�ʭs�쒿nP��a�ǿN���2��ֈ����H�
����ֈ��2��x   x   �$��t�����ɭs��tH�x6"��"��ҾO����.!��/!������S�Ҿ�"�w6"��tH���s���u����$���$տ�濧��!w��!w��������$տx   x   \����؋���m��2F�x6"��F���ԾsD���m��7:��P:��0:���m��cD����Ծ�F�z6"��2F���m��؋�\���g8���3ſ�bҿY�ڿD�ݿR�ڿcҿ�3ſe8��x   x   H�����b�L�?�����"���Ծ_����ꔾh��o�u�j�u�h���ꔾg�����Ծ�"����O�?���b�F������٤�>뱿�?���������?��=뱿�٤���x   x   �jS�l95�t��1����ҾsD���ꔾ�|��oGo�!h�tGo��|���ꔾoD���Ҿ1���v��h95��jS��q��䆿D$�����ˤ��г��ˤ�����C$���䆿�q�x   x    �'�
��Z�
7;O�m��h��oGo�
�c��c�{Go�h���m��M
7;Z���'�'�ݩ@�^�X�؉n�[B��|���������}���^B��։n�`�X��@�x   x   P5��c��ƾb������7:��o�u�!h��c�	!h�r�u�2:������O���ƾ�c�U5�i����+�P>��BN�u�Z�	vb�%e�vb�t�Z��BN�P>���+�l��x   x   (�׾BR��&���.!��P:��j�u�tGo�{Go�r�u�N:��-!���&��JR��)�׾���MU�>��>�#��.��6��:��:���6��.�:�#�B��LU����x   x   Bط�&���,���[��/!��0:��h���|��h��2:��-!���[��,��*���:ط��`ɾ�ܾ!��(���
�������h��������
�(�1��دܾ�`ɾx   x   `5���<��,��������m���ꔾ�ꔾ�m�������,���<��\5�����挻��@Ǿ�\Ӿ��޾~�辜�������辺�޾�\Ӿ�@Ǿ،�����x   x   f5��$���&��Z��ScD��g���oD��MO��&��*���\5��`
��)t��[@��������R����	þ��žQ�ƾ��ž�	þM���������`@��t��f
��x   x   @ط�?R���ƾ7;�Ҿ��Ծ��Ծ�Ҿ
7;�ƾJR��:ط����)t���\��褾�̣�ɯ��%��5����$���$��;���%%��Ư���̣�	褾�\��t�����x   x   2�׾�c�&Z�,����"��F��"�1���Z��c�)�׾�`ɾ挻�[@��褾����rp����$A�������-������.A����sp�������社a@��ڌ���`ɾx   x   R5���z�����w6"�z6"����v����U5�����ܾ�@Ǿ����̣�rp��������(��#�z��z�2��������wp���̣�����@Ǿ�ܾ���x   x   %�'�h95�S�?��2F��tH��2F�O�?�h95�'�'�i��MU�!���\Ӿ���ɯ���������v��wk���g��wk��v������ǯ������\Ӿ&��OU�d��x   x   �jS���b���m�ʭs���s���m���b��jS�ݩ@���+�>��(���޾R���%��$A��(���wk���a��a��wk�2��,A��%��W�����޾(�>����+�ک@�x   x   F����؋���쒿���؋�F����q�^�X�P>�>�#���
�~���	þ5�������#�z���g��a���g��z�����<����	þ��辷�
�=�#�P>�b�X��q�x   x   \���t���lP��nP��u���\������䆿؉n��BN��.�������ž�$���-���z��wk��wk��z��-���$����ž�����.��BN�։n��䆿��x   x   �$��e�ǿ;Jʿa�ǿ�$��g8���٤�D$��[B��u�Z��6�������Q�ƾ�$������2���v�2�������$��L�ƾ�������6�t�Z�`B��C$���٤�g8��x   x   O��5}�6}�N���$տ�3ſ>뱿���|���	vb��:��h������ž;���.A��������,A��<�����ž��� i��:�vb�}������=뱿�3ſ�$տx   x   ( �x��( ��2�����bҿ�?��ˤ�����%e��:�������	þ%%���������%���	þ������:�%e����ˤ���?��cҿ���2��x   x   %��'��r�
�ֈ����Y�ڿ���г�����vb���6������M���Ư��sp��wp��ǯ��W���������6�vb����ҳ�����O�ڿ���و�p�
�x   x   ���uw� h����!w��D�ݿ���ˤ��}���t�Z��.���
���޾����̣������̣������޾��
��.�t�Z�}���ˤ�����D�ݿ!w����� h�uw�x   x   �:#�o��bj�H�
�!w��R�ڿ�?�����^B���BN�:�#�(��\Ӿ���	褾�社����\Ӿ(�=�#��BN�`B������?��O�ڿ!w��I�
�aj�n���:#�x   x   ��'�!�`j�������cҿ=뱿C$��։n�P>�B��1���@Ǿ`@���\��a@���@Ǿ&��>��P>�։n�C$��=뱿cҿ�����aj�!���'� *�x   x   ��'�o��h�ֈ��濇3ſ�٤��䆿`�X���+�LU�دܾ،��t��t��ڌ���ܾOU���+�b�X��䆿�٤��3ſ��و� h�n����'�},�},�x   x   �:#�sw�s�
��2���$տe8�����q��@�l������`ɾ���f
������`ɾ���d��ک@��q���g8���$տ�2��p�
�uw��:#� *�},�*�x   x   �L� ��,�׿R������H���{�U�E++�J���۾�o���l��Rz���l���o����۾J�E++�~�U�I�������R��-�׿��L�%��pb�g�nb�&��x   x    ���ڿ2���Ӥ�(-����b�N7�9��<꾈O��hj��<:��=:��lj���O���<�9�M7���b�'-���Ӥ�2����ڿ����p�
�ǂ�Ȃ�r�
���x   x   ,�׿2��Y�����L3k�L�?�_��י��LjȾ�è�`J��q-��[J���è�QjȾݙ��Z��M�?�B3k�����W�2��1�׿�쿯���و�;K�׈�������x   x   R���Ӥ�����gn�+D���������ξT﫾wS��0-��2-��yS��N﫾��ξ������(D�on������Ӥ�R��>�Ͽۗ࿏�쿨���򿍫�ח�@�Ͽx   x   ����(-��L3k�+D��� ��"�7.Ӿg������� ������ ������ g��;.Ӿ�"��� �*D�P3k�'-������M����¿��ϿF�׿O�ڿH�׿��Ͽ�¿N���x   x   H�����b�L�?�����"���Ծ_����ꔾh��o�u�j�u�h���ꔾg�����Ծ�"����O�?���b�F������٤�>뱿�?���������?��=뱿�٤���x   x   {�U�N7�_�����7.Ӿ_���픾m+��u@n�G�f��@n�r+��픾d���?.Ӿ���Y��L7�x�U�c]t����+���b���γ���ʦ�ҳ��_���)������^]t�x   x   E++�9�י����ξg���ꔾm+��	�k�x�_�u�_���k�o+���ꔾg����ξљ��9�C++���D��]�7t��c������s���s������c��7t��]���D�x   x   J��<�LjȾT﫾����h��u@n�x�_�|�Z�s�_�@n�h������V﫾NjȾ�<�J�i���L1���D�XqU�vb�z�j�[�m�z�j�vb�YqU���D��L1�l��x   x   ��۾�O���è�wS��� ��o�u�G�f�u�_�s�_�I�f�g�u�� ��{S���è��O����۾������������*��6�R�>�B`C�H`C�U�>��6���*����������x   x   �o��hj��`J��0-�����j�u��@n���k�@n�g�u����.-��fJ��aj���o����˾�_�ow��P�����6���������6���T��lw���_���˾x   x   �l��<:��q-��2-��� ��h��r+��o+��h��� ��.-��n-��;:���l������~���s˾D�ھx����������r�w�~����������D�ھ�s˾~������x   x   Rz��=:��[J��yS�������ꔾ픾�ꔾ����{S��fJ��;:��Lz��^@��i�������P��J���Rbƾ��̾ �о;	Ҿ/�о��̾SbƾW����P�����^���Z@��x   x   �l��lj���è�N﫾 g��g���d���g��V﫾�è�aj���l��^@���G�������?������@���N��|��������%|���M��F���ǯ���?�������G��T@��x   x   �o���O��QjȾ��ξ;.Ӿ��Ծ?.Ӿ��ξNjȾ�O���o������i��������H��np����q|��(����s���`���s��#���k|����wp���H������]�������x   x   ��۾�<�ݙ������"��"����љ���<꾞�۾��˾~������?��np��vȍ��8������J��u|��u|�J������8��|ȍ�sp���?�����~����˾x   x   J�9�Z������� ����Y��9�J������_⾇s˾�P���������8���,{��m���e�=@c���e��m��,{��8����Ư���P���s˾�_⾐���x   x   E++�M7�M�?�(D�*D�O�?�L7�C++�i�����ow��D�ھJ���@���q|�������m�ve^�>�V�L�V�}e^��m�����r|��F���M���:�ھhw�����l��x   x   ~�U���b�B3k�on�P3k���b�x�U���D��L1����P��x��RbƾN��(���J���e�>�V���Q�7�V���e��I�$���N��Sbƾ���Q�����L1���D�x   x   I���'-����������'-��F���c]t��]���D���*���������̾|���s���u|�=@c�L�V�7�V�N@c�}u|��s��|����̾��������*���D��]�d]t�x   x   �����Ӥ�W��Ӥ� ��������7t�XqU��6��6����� �о����`���u|���e�}e^���e�}u|��`�����)�о�����6���6�VqU�7t�!�����x   x   R��2��2��R��M����٤�+����c��vb�R�>���r�;	Ҿ����s��J��m��m��I��s�����H	Ҿt���U�>�vb��c��,����٤�P���x   x   -�׿��ڿ1�׿>�Ͽ�¿>뱿b������z�j�B`C����w�/�о%|��#��������,{�����$���|��)�оt����G`C�z�j����b���<뱿�¿@�Ͽx   x   ������ۗ࿰�Ͽ�?��γ���s��[�m�H`C���~�����̾�M��k|���8���8��r|��N����̾������G`C�P�m��s��г���?����Ͽؗ���x   x   �L����������F�׿����ʦ��s��z�j�U�>��6�����SbƾF�����|ȍ���F���Sbƾ�����6�U�>�z�j��s���ʦ����F�׿��쿯�����x   x   %��p�
�و����O�ڿ���ҳ�����vb��6������W���ǯ��wp��sp��Ư��M����������6�vb����г�����Y�ڿ���ֈ�r�
�'��x   x   pb�ǂ�;K����H�׿�?��_����c��YqU���*�T��D�ھ�P���?���H���?���P��:�ھQ����*�VqU��c��b����?��F�׿���<K�Ȃ�ob�&g�x   x   g�Ȃ�׈���쿯�Ͽ=뱿)���7t���D���lw���s˾���������������s˾hw������D�7t�,���<뱿��Ͽ���ֈ�Ȃ�	g�͈�͈�x   x   nb�r�
�����ח��¿�٤�����]��L1�����_�~��^����G��]���~���_⾬���L1��]�!����٤��¿ؗ࿯���r�
�ob�͈���͈�x   x   &������@�ϿN�����^]t���D�l��������˾����Z@��T@��������˾����l����D�d]t���P���@�Ͽ����'��&g�͈�͈�&g�x   x   r�࿷xʿN�� 𘿬q���jS�E++�k[	���ݾ~l���מ�K���O����מ�|l����ݾh[	�H++��jS��q��!�K���xʿr����( ���	��' ���x   x   �xʿd\���؜��L����]�l95�9����q���ʠ��*w��eΌ�,w��Ϡ��u������9�g95���]��L���؜�d\���xʿ~�ݿ���2���u���2����}�ݿx   x   N���؜������:c�j�;�t��י���ɾ,��K钾�j���j��I钾
,���ɾԙ��v��o�;��:c������؜�N���Mſ�6տؗ�����՗��6տ�Mſx   x    ��L���:c��=�V��1�����ξ$�U����f�� ����f��U���'���ξ=���U���=��:c��L��!��^��ga��v�ǿ��Ͽcҿ��Ͽv�ǿga���^��x   x   �q����]�j�;�V���	 ��Ҿg���s������W[v�V[v������s��g���Ҿ|	 �U��h�;���]��q���m��cˠ�nz��N����?���?��M���oz��aˠ��m��x   x   �jS�l95�t��1����ҾsD���ꔾ�|��oGo�!h�tGo��|���ꔾoD���Ҿ1���v��h95��jS��q��䆿D$�����ˤ��г��ˤ�����C$���䆿�q�x   x   E++�9�י����ξg���ꔾm+��	�k�x�_�u�_���k�o+���ꔾg����ξљ��9�C++���D��]�7t��c������s���s������c��7t��]���D�x   x   k[	���뾜ɾ$��s���|��	�k�]��X�]��k��|���s��'��ɾ��h[	�u4�t!3�{�F�w�W�%e�O�m�afp�P�m�%e�t�W�z�F�x!3�v4�x   x   ��ݾq���,��U�������oGo�x�_��X��X�|�_�oGo�����V���	,��t�����ݾJb���N�0���c.��:�F`C�`�G�_�G�G`C��:��c.�4���N�Hb��x   x   ~l��ʠ��K钾�f��W[v�!h�u�_�]�|�_�!h�T[v��f��K钾Ơ���l��#�;�&澃��x�������=#��%��=#������~x�����&��;x   x   �מ�*w���j�� ���V[v�tGo���k��k�oGo�T[v������j��(w���מ�R��Ӄ����ξ�߾�𾉊������3��3�����������߾��ξك��R��x   x   J���eΌ��j���f�������|��o+���|�������f���j��jΌ�O���r[��Jj�����)k���	þ��̾%5Ծ# پ{�ھ( پ%5Ծ��̾�	þ'k��,���Vj��e[��x   x   O���,w��I钾U����s���ꔾ�ꔾ�s��V���K钾(w��O������i����V������%%��N��d߭�(K��������'K��d߭�N��%�������V��t������x   x   �מ�Ϡ��
,��'�g��oD��g��'�	,��Ơ���מ�r[��i������x����v|���W��6O������Q�����BO���W��r|�����x����o���f[��x   x   |l��u����ɾ��ξ�Ҿ�Ҿ��ξ�ɾt����l��R��Jj���V���x�����9��\����b��� ���~�0�~�� ���b��b����8������x���V��[j��R��x   x   ��ݾ���ԙ��=���|	 �1���љ���뾤�ݾ#�;Ӄ�����������9��,$}��p�x"g���a��*`���a�w"g��p�*$}��8��������-���΃��#�;x   x   h[	�9�v��U��U��v��9�h[	�Jb���&澤�ξ)k��%%��v|��\����p�6�^�ۨS��N�~N��S�/�^��p�b���k|��%%��$k����ξ�&�Vb��x   x   H++�g95�o�;��=�h�;�h95�C++�u4��N�����߾�	þN���W���b��x"g�ۨS��H��CD��H��S��"g��b���W���M���	þ�߾����N�n4�x   x   �jS���]��:c��:c���]��jS���D�t!3�0��x��𾤗̾d߭�6O��� ����a��N��CD��CD��N���a�� ��8O��d߭���̾��x�4��x!3���D�x   x   �q���L�������L���q���q��]�{�F��c.��������%5Ծ)K������~��*`�~N��H��N��*`�2�~����*K��%5Ծ~�������c.�y�F��]��q�x   x   !𘿽؜��؜�!𘿺m���䆿7t�w�W��:������# پ����Q��0�~���a��S��S���a�2�~��Q�����  پ������:��W�7t��䆿�m��x   x   K��d\��N���^��cˠ�D$���c��%e�F`C��=#��3�{�ھ������� ��w"g�/�^��"g�� ��������t�ھ�3��=#�H`C�%e��c��@$��cˠ��^��x   x   �xʿ�xʿ�Mſga��nz��������O�m�`�G��%��3�( پ'K��BO���b���p��p��b��8O��*K��  پ�3��%�_�G�[�m�������nz��ba���Mſx   x   r��~�ݿ�6տv�ǿN���ˤ���s��afp�_�G��=#����%5Ծd߭��W��b���*$}�b����W��d߭�%5Ծ����=#�_�G�afp��s��ˤ��N���v�ǿ�6տ~�ݿx   x   ����ؗ࿳�Ͽ�?��г���s��P�m�G`C���������̾N��r|���8���8��k|���M����̾~�����H`C�[�m��s��γ���?����Ͽۗ�����x   x   ( ��2����cҿ�?��ˤ�����%e��:�������	þ%���������%%���	þ������:�%e����ˤ���?���bҿ���2��( �x��x   x   ���u���濶�ϿM�������c��t�W��c.�~x��߾'k�������x���x������$k���߾�x��c.��W��c�����N�����Ͽ���u����i�k�x   x   	���2��՗�v�ǿoz��C$��7t�{�F�4�������ξ,����V�����V��-�����ξ���4��y�F�7t�@$��nz��v�ǿۗ��2�������c�
����x   x   ' ����6տga��aˠ��䆿�]�x!3��N��&�ك��Vj��t���o���[j��΃���&��N�x!3��]��䆿cˠ�ba���6տ��( �i�c�
�b�
�j�x   x   ��}�ݿ�Mſ�^���m���q���D�v4�Hb���;R��e[�����f[��R��#�;Vb��n4���D��q��m���^���Mſ~�ݿ��x��k����j�z��x   x   ������2ُ�ou�ڍL� �'�J���ݾ'v���$��߭��Q���ݭ���$��(v����ݾJ�%�'��L�ju�/ُ��������xʿ-�׿O�࿛{�Q��,�׿�xʿx   x   ���٪��\7{�oT�3�/�
���<�q���Q��⩏�[��\��穏�V��u����<���0�/�lT�W7{�ݪ�����i����Mſ@�Ͽ�$տ�$տ@�Ͽ�Mſk���x   x   2ُ�\7{�0�V�:�3���Z�LjȾ,��Fϑ�����mG������?ϑ�	,��MjȾZ���;�3�)�V�[7{�1ُ�����xׯ�ba���¿�3ſ�¿ea��vׯ�����x   x   ou�oT�:�3��$�w ��
7;T﫾U���5Ճ��x��x�4Ճ�^���N﫾7;l ���$�:�3�wT�pu�È�������nz��<뱿=뱿nz���󤿫��ƈ��x   x   ڍL�3�/���w ����ξO��������Pwr���k�Uwr���������P��ξ} ����0�/�ݍL��Ki��!��ԍ��䖿���b�������䖿ԍ��!���Ki�x   x    �'�
��Z�
7;O�m��h��oGo�
�c��c�{Go�h���m��M
7;Z���'�'�ݩ@�^�X�؉n�[B��|���������}���^B��։n�`�X��@�x   x   J��<�LjȾT﫾����h��u@n�x�_�|�Z�s�_�@n�h������V﫾NjȾ�<�J�i���L1���D�XqU�vb�z�j�[�m�z�j�vb�YqU���D��L1�l��x   x   ��ݾq���,��U�������oGo�x�_��X��X�|�_�oGo�����V���	,��t�����ݾJb���N�0���c.��:�F`C�`�G�_�G�G`C��:��c.�4���N�Hb��x   x   'v��Q��Fϑ�5Ճ�Pwr�
�c�|�Z��X�g�Z��c�^wr�9Ճ�Bϑ�T��$v��y�ξUy�ۅ ���� i�����%���&��%���� i����ޅ �Ly�v�ξx   x   �$��⩏������x���k��c�s�_�|�_��c���k��x�����詏��$���Ȭ�'���о��⾓��v��3�*��1���3�t��������о'���Ȭ�x   x   ߭��[��mG���x�Uwr�{Go�@n�oGo�^wr��x�tG��X��ޭ��T���,�������)빾��ž,�о پj�޾fz�i�޾  پ)�о��ž#빾����3���Y���x   x   Q���\������4Ճ�����h��h������9Ճ�����X��K���^7����������/���!|�� K������ַ��ַ����+K��|��<������{����Z7��x   x   ݭ��穏�?ϑ�^��������m������V���Bϑ�詏�ޭ��^7��O���P㋾�+��$A��"���1O������1������,������8O��$���,A���+��B㋾Q���_7��x   x   �$��V��	,��N﫾PMV﫾	,��T���$��T�����P㋾巇��������c��Ӏ�%���n���l���-���Ӏ��b���������𷇾B㋾��Y���x   x   (v��v���MjȾ7;��ξ
7;NjȾt���$v���Ȭ�,�������+������,{��p�+�g� }b�W_�qQ^�W_��|b�$�g��p��,{�����+����.����Ȭ�x   x   ��ݾ�<�Z�l ��} ��Z��<꾤�ݾy�ξ'���������$A�������p�{�_��RS�MVK�
fG��eG�MVK��RS�i�_��p�����.A��
�������'��x�ξx   x   J������$�����J�Jb��Uy��о)빾/���"���c��+�g��RS���D��<��'9��<���D��RS�$�g��b��#���;���빾�оOy�Bb��x   x   %�'�0�/�;�3�:�3�0�/�'�'�i���N�ۅ ������ž!|��1O��Ӏ� }b�MVK��<�fm4�ym4��<�KVK��|b�Ӏ�BO��%|����ž���څ ��N�l��x   x   �L�lT�)�V�wT�ݍL�ݩ@��L1�0��������,�о K������%���W_�
fG��'9�ym4��'9��eG�W_��������'K��.�о��󾰹�2�� M1�ީ@�x   x   ju�W7{�[7{�pu��Ki�^�X���D��c.� i�v� پ���1��n���qQ^��eG��<��<��eG�`Q^�i���0�����( پw��h��c.���D�d�X��Ki�x   x   /ُ�ݪ��1ُ�È���!��؉n�XqU��:�����3�j�޾�ַ�����l���W_�MVK���D�KVK�W_�i��������ַ�i�޾�3�����:�YqU�׉n��!��ň��x   x   �������������ԍ�[B��vb�F`C��%�*��fz��ַ�,��-����|b��RS��RS��|b����0���ַ�uz�1���%�B`C�	vb�_B��ԍ��������x   x   ���i���xׯ��󤿊䖿|���z�j�`�G���&�1��i�޾�������Ӏ�$�g�i�_�$�g�Ӏ��������i�޾1����&�`�G�z�j�|����䖿��xׯ�i���x   x   �xʿ�Mſba��nz��������[�m�_�G��%��3�  پ+K��8O���b���p��p��b��BO��'K��( پ�3��%�`�G�O�m�������nz��ga���Mſ�xʿx   x   -�׿@�Ͽ�¿<뱿b������z�j�G`C����t�)�о|��$��������,{�����#���%|��.�оw����B`C�z�j����b���>뱿�¿>�Ͽ1�׿��ڿx   x   O���$տ�3ſ=뱿���}���vb��:� i������ž<���,A��������.A��;�����ž����h��:�	vb�|������>뱿�3ſ�$տN��6}�5}�x   x   �{��$տ�¿nz���䖿^B��YqU��c.�������#빾����+��𷇾�+��
���빾��⾰���c.�YqU�_B���䖿nz���¿�$տ�{�������x   x   Q��@�Ͽea����ԍ�։n���D�4��ޅ ��о����{��B㋾B㋾�������оڅ �2����D�։n�ԍ���ga��>�ϿN����m��l����x   x   ,�׿�Mſvׯ�����!��`�X��L1��N�Ly�'��3�����Q�����.���'��Oy��N� M1�d�X��!�����xׯ��Mſ1�׿6}���l����2}�x   x   �xʿk�������ƈ���Ki��@�l��Hb��v�ξ�Ȭ�Y���Z7��_7��Y����Ȭ�x�ξBb��l��ީ@��Ki�ň������i����xʿ��ڿ5}�����2}濐�ڿx   x   �p���!���d�a�A���!�P5���۾~l���$�����9���8�������$��l����۾O5���!�`�A���d��!���p�����K��R���$���$��R��M�����x   x   �!��=cg�xF��;'����c澈O��ʠ��⩏�/郾���0郾婏�Ǡ���O���c澑��;'�xF�Ccg��!����������^��P���g8��O����^���������x   x   �d�xF�00)�J.��C��ƾ�è�K钾����P1{�J1{�����H钾�è��ƾ�C�N.�/0)�xF�w�d�b���������cˠ��٤��٤�cˠ�������a���x   x   a�A��;'�J.����ʾb��wS���f���x� �q��x��f��zS��^��ʾx��I.��;'�^�A�L\��;u��p��ԍ�@$��,���C$��ԍ��p���;u�L\�x   x   ��!����C�ʾ5������� ��W[v���k���k�T[v�� ������5��ʾ�C��}�!���8��9O�g�c��~t�_B���c���c��`B���~t�f�c��9O���8�x   x   P5��c��ƾb������7:��o�u�!h��c�	!h�r�u�2:������O���ƾ�c�U5�i����+�P>��BN�u�Z�	vb�%e�vb�t�Z��BN�P>���+�l��x   x   ��۾�O���è�wS��� ��o�u�G�f�u�_�s�_�I�f�g�u�� ��{S���è��O����۾������������*��6�R�>�B`C�H`C�U�>��6���*����������x   x   ~l��ʠ��K钾�f��W[v�!h�u�_�]�|�_�!h�T[v��f��K钾Ơ���l��#�;�&澃��x�������=#��%��=#������~x�����&��;x   x   �$��⩏������x���k��c�s�_�|�_��c���k��x�����詏��$���Ȭ�'���о��⾓��v��3�*��1���3�t��������о'���Ȭ�x   x   ���/郾P1{� �q���k�	!h�I�f�!h���k��q�E1{�.郾��������0��ۘ���u��B�ƾ<	Ҿ��ھkzྀm�uz�t�ھH	ҾL�ƾ�u��瘭��0������x   x   9������J1{��x�T[v�r�u�g�u�T[v��x�E1{����:����^���\���l��-���$���������ַ��T���T���ַ��������$��-���l���\���^��x   x   8���0郾�����f��� ��2:��� ���f������.郾:��������.����������s�����=��������������0������s����������.������x   x   ���婏�H钾zS����������{S��K钾詏�����^�����׀������9��J�� ��)����:������ȕ���:������ ���I�2������ـ������^��x   x   �$��Ǡ���è�^��5��O���è�Ơ���$�������\���.�������v�(�m�w"g��|b�q�_���]��[]���]���_��|b��"g��m��v������.���\������x   x   l���O���ƾʾʾ�ƾ�O���l���Ȭ��0���l�����9��(�m�7�^��RS���J��UE���B���B��UE���J��RS�/�^��m�2������l���0���Ȭ�x   x   ��۾�c澪C�x�ﾞC��c澞�۾#�;'��ۘ��-������J�x"g��RS��D�9,9��2�Ι0���2�B,9��D��RS�w"g�J�����-��옭�'���;x   x   O5���N.�I.���U5������&��о�u���$���s��� ���|b���J�9,9� u-��'��'��t-�B,9���J��|b�� ���s���$���u���о�&澉���x   x   ��!��;'�/0)��;'�}�!�i�����������B�ƾ������)���q�_��UE��2��'�h�#���'���2��UE���_�-���������Q�ƾ��⾅�����f��x   x   `�A�xF�xF�^�A���8���+����x����<	Ҿ���=���:����]���B�Ι0��'���'�ߙ0���B���]��:��,�����;	Ҿ���x�����+���8�x   x   ��d�Ccg�w�d�L\��9O�P>���*����v���ھ�ַ����������[]���B���2��t-���2���B��[]�ƕ�������ַ�{�ھr������*�P>��9O�L\�x   x   �!���!��b����;u�g�c��BN��6����3�kz��T������ȕ����]��UE�B,9�B,9��UE���]�ƕ�������T��fzྱ3����6��BN�b�c��;u�d���x   x   �p���������p���~t�u�Z�R�>��=#�*���m��T�������:����_���J��D���J���_��:�������T���m�*���=#�R�>�u�Z��~t��p��������x   x   ����������ԍ�_B��	vb�B`C��%�1��uz��ַ�0������|b��RS��RS��|b�-���,���ַ�fz�*���%�F`C�vb�[B��ԍ�����������x   x   K���^��cˠ�@$���c��%e�H`C��=#��3�t�ھ������� ���"g�/�^�w"g�� ��������{�ھ�3��=#�F`C�%e��c��D$��cˠ��^��N��d\��x   x   R��P����٤�,����c��vb�U�>���t�H	Ҿ����s���I��m��m�J��s�����;	Ҿr���R�>�vb��c��+����٤�M���R��2��2��x   x   �$��g8���٤�C$��`B��t�Z��6�������L�ƾ�$������2���v�2�������$��Q�ƾ�������6�u�Z�[B��D$���٤�g8���$��a�ǿ;Jʿe�ǿx   x   �$��O���cˠ�ԍ��~t��BN���*�~x�����u��-����������������-���u����⾀x���*��BN��~t�ԍ�cˠ�M����$���Eʿ!�Ͽ"�Ͽ�Eʿx   x   R���^������p��f�c�P>�������о瘭��l���.��ـ���.���l��옭��о�����P>�b�c��p������^��R��a�ǿ!�Ͽ�=ҿ!�Ͽ`�ǿx   x   M����������;u��9O���+�����&�'���0���\���������\���0��'���&澫����+��9O��;u��������N��2��;Jʿ"�Ͽ!�Ͽ=Jʿ2��x   x   ������a���L\���8�l�������;�Ȭ������^����^�������Ȭ��;����f����8�L\�d���������d\��2��e�ǿ�Eʿ`�ǿ2��f\��x   x   �Im�e�P���3�!���u �(�׾�o���מ�߭��9���vG��>���᭍��מ��o��(�׾�u �#����3�_�P��Im��!��/ُ�!�����\������� �/ُ��!��x   x   e�P�6��Q�H��B��BR��hj��*w��[��������W��1w��jj��GR��F��A���Q�6�g�P��_j�d���ň���m�������m��È��f����_j�x   x   ��3��Q�_+�C�-Wľ&��`J���j��mG��J1{�qG���j��WJ��&��&WľE�d+��Q���3���K� �a��;u��!���䆿!����䆿�!���;u� �a���K�x   x   !��H��C�Cƾ�����0-�� ����x��x�����2-�������Hƾ<�H��"����-���A��`T�b�c�׉n�7t�7t�։n�]�c��`T���A���-�x   x   �u �B��-Wľ�������.!�����V[v�Uwr�T[v����.!���������+WľI���u �����#��X4���B��BN�YqU��W�VqU��BN���B��X4���#���x   x   (�׾BR��&���.!��P:��j�u�tGo�{Go�r�u�N:��-!���&��JR��)�׾���MU�>��>�#��.��6��:��:���6��.�:�#�B��LU����x   x   �o��hj��`J��0-�����j�u��@n���k�@n�g�u����.-��fJ��aj���o����˾�_�ow��P�����6���������6���T��lw���_���˾x   x   �מ�*w���j�� ���V[v�tGo���k��k�oGo�T[v������j��(w���מ�R��Ӄ����ξ�߾�𾉊������3��3�����������߾��ξك��R��x   x   ߭��[��mG���x�Uwr�{Go�@n�oGo�^wr��x�tG��X��ޭ��T���,�������)빾��ž,�о پj�޾fz�i�޾  پ)�о��ž#빾����3���Y���x   x   9������J1{��x�T[v�r�u�g�u�T[v��x�E1{����:����^���\���l��-���$���������ַ��T���T���ַ��������$��-���l���\���^��x   x   vG�����qG���������N:���������tG�����xG���5������%��� ���-���`���Q�����������h�����������Q���`���-����%��������5��x   x   >���W���j��2-��.!��-!��.-���j��X��:����5���v~��{�B�z��z�yu|�$�~�m���Ǖ���%���%��ƕ��i���2�~�}u|��z�=�z��{��v~��5��x   x   ᭍�1w��WJ�������fJ��(w��ޭ���^�������{�	�r��wk���e���a�W_���]��(]��\��(]���]�W_���a���e��wk���r��{������^��x   x   �מ�jj��&����������&��aj���מ�T����\��%���B�z��wk�oe^�ܨS�OVK��UE�|A���?���?��{A��UE�KVK��S�}e^��wk�A�z�����\��R���x   x   �o��GR��&WľHƾ+WľJR���o��R��,����l�� ���z���e�ܨS���D�<,9�`1�N/,���*�[/,�M1�B,9���D��S���e��z����l��(���R��x   x   (�׾F��E�<�I��)�׾��˾Ӄ������-���-��yu|���a�OVK�<,9���+���"�������"�}�+�B,9�MVK���a��u|��-��-������у���˾x   x   �u �A��d+�H���u ����_⾤�ξ)빾�$���`��$�~�W_��UE�`1���"������������"�M1��UE�W_�0�~��`���$��빾��ξ�_⾒��x   x   #���Q��Q�"����MU�ow���߾��ž����Q��m�����]�|A�N/,�����������?/,��{A���]�l����Q�������ž�߾gw��PU���x   x   ��3�6���3���-���#�>��P����,�о�������Ǖ���(]���?���*����������*���?��(]�ȕ��������� �о��R��C����#���-�x   x   _�P�g�P���K���A��X4�?�#������� پ�ַ������%���\���?�[/,���"���"�?/,���?�
�\��%�������ַ�# پ������=�#��X4���A���K�x   x   �Im��_j� �a��`T���B��.��6����j�޾�T���h���%���(]��{A�N1�}�+�M1��{A��(]��%���h���T��j�޾����6��.���B��`T� �a��_j�x   x   �!��d����;u�b�c��BN��6����3�fz��T������ƕ����]��UE�B,9�B,9��UE���]�ȕ�������T��kzྫ3����6��BN�g�c��;u�b����!��x   x   /ُ�ň���!��׉n�YqU��:�����3�i�޾�ַ�����i���W_�KVK���D�MVK�W_�l��������ַ�j�޾�3�����:�XqU�؉n��!��È��1ُ�ݪ��x   x   !𘿹m���䆿7t��W��:������  پ����Q��2�~���a��S��S���a�0�~��Q�����# پ������:�w�W�7t��䆿�m��!𘿻؜��؜�x   x   ������!���7t�VqU���6��6�����)�о����`��}u|���e�}e^���e��u|��`����� �о�����6��6�XqU�7t�����������Ӥ�W��Ӥ�x   x   \������䆿׉n��BN��.�������ž�$���-���z��wk��wk��z��-���$����ž�����.��BN�؉n��䆿��\���u���nP��lP��t���x   x   �����m���!��]�c���B�:�#�T���߾#빾-����=�z���r�A�z���-��빾�߾R��=�#���B�g�c��!���m������u�������滱�����v���x   x    �È���;u��`T��X4�B��lw����ξ�����l��%����{��{�����l��������ξgw��C���X4��`T��;u�È��!��Ӥ�nP��滱�仱�lP���Ӥ�x   x   /ُ�f��� �a���A���#�LU��_�ك��3����\�������v~������\��(���у���_�PU���#���A� �a�b���1ُ��؜�W�lP������lP��Y��؜�x   x   �!���_j���K���-��������˾R��Y����^���5���5���^��R���R���˾�������-���K��_j��!��ݪ���؜��Ӥ�t���v����Ӥ��؜�ߪ��x   x   O�:�$��R��$��F`ӾBط��l��K���Q���8���>���L���M����l��6ط�X`Ӿ�$���R�$�G�:�_�P���d�ju��q��I���F����q��nu�y�d�^�P�x   x   $���w����پ}r��&���<:��eΌ�\��0郾W��fΌ�@:��0����r����پw�����$��]8���K�L\��Ki��q�d]t��q��Ki�L\���K��]8�x   x   �R�w��2�۾H���̮��,��q-���j�����������j��j-��,��Ǯ��J���J�۾w���R��> ���1���A��9O�d�X��]��]�b�X��9O���A���1��> �x   x   �$����پH�������=���[��2-���f��4Ճ��f��2-���[���=�����C�����پ�$����	������'��X4�P>���D�y�F���D�P>��X4���'������	�x   x   F`Ӿ}r��̮���=����/!��� ����������� ��.!�����=��®���r��Q`Ӿ���x�!���5�=�#���*��c.��c.���*�=�#��5� ��w����x   x   Bط�&���,���[��/!��0:��h���|��h��2:��-!���[��,��*���:ط��`ɾ�ܾ!��(���
�������h��������
�(�1��دܾ�`ɾx   x   �l��<:��q-��2-��� ��h��r+��o+��h��� ��.-��n-��;:���l������~���s˾D�ھx����������r�w�~����������D�ھ�s˾~������x   x   K���eΌ��j���f�������|��o+���|�������f���j��jΌ�O���r[��Jj�����)k���	þ��̾%5Ծ# پ{�ھ( پ%5Ծ��̾�	þ'k��,���Vj��e[��x   x   Q���\������4Ճ�����h��h������9Ճ�����X��K���^7����������/���!|�� K������ַ��ַ����+K��|��<������{����Z7��x   x   8���0郾�����f��� ��2:��� ���f������.郾:��������.����������s�����=��������������0������s����������.������x   x   >���W���j��2-��.!��-!��.-���j��X��:����5���v~��{�B�z��z�yu|�$�~�m���Ǖ���%���%��ƕ��i���2�~�}u|��z�=�z��{��v~��5��x   x   L���fΌ�j-���[�����[��n-��jΌ�K�����v~���u���m���g�<@c��*`�|Q^��[]��\���\�
�\��[]�`Q^��*`�N@c���g���m���u��v~��x   x   M���@:��,���=���=��,��;:��O���^7������{���m�
�a�I�V��N��eG���B���?��'>��'>���?���B��eG��N�7�V��a���m�!�{����[7��x   x   �l��0���Ǯ�����®��*����l��r[�����.��B�z���g�I�V��H��<���2�M/,�O(�'�O(�?/,���2��<��H�L�V���g�E�z��.����p[��x   x   6ط��r��J���C����r��:ط�����Jj���������z�<@c��N��<��t-���"�Q>������j>���"��t-��<�}N�=@c�#�z�������Hj������x   x   X`Ӿ��پJ�۾��پQ`Ӿ�`ɾ~������������yu|��*`��eG���2���"���������}�������"���2��eG��*`��u|��������'���~���`ɾx   x   �$��w��w���$������ܾ�s˾)k��/����s��$�~�|Q^���B�M/,�Q>�����D
��D
����j>�[/,���B�qQ^��~��s��5���2k���s˾ܾ߯���x   x   �R�����R���	�x�!��D�ھ�	þ!|�����m����[]���?�O(�������D
�����O(���?��[]�n������|���	þA�ھ+��v��	�x   x   $�$��> ����!��(�x�辤�̾ K��=��Ǖ���\��'>�'���}�������,'��'>��\�����1��(K����̾~��(�������> �x   x   G�:��]8���1���'��5���
�����%5Ծ��������%����\��'>�O(�j>����j>�O(��'>���\��%���������%5Ծ������
��5���'���1��]8�x   x   _�P���K���A��X4�=�#�������# پ�ַ������%��
�\���?�?/,���"���"�[/,���?��\��%�������ַ� پ������>�#��X4���A���K�g�P�x   x   ��d�L\��9O�P>���*����r�{�ھ�ַ�����ƕ���[]���B���2��t-���2���B��[]����������ַ���ھv������*�P>��9O�L\�w�d�Ccg�x   x   ju��Ki�d�X���D��c.��h�w�( پ���0��i���`Q^��eG��<��<��eG�qQ^�n���1����� پv� i��c.���D�^�X��Ki�pu�[7{�W7{�x   x   �q���q��]�y�F��c.����~���%5Ծ+K�����2�~��*`��N��H�}N��*`��~����(K��%5Ծ��������c.�{�F��]��q��q���L�������L��x   x   I���d]t��]���D���*���������̾|���s��}u|�N@c�7�V�L�V�=@c��u|��s��|����̾��������*���D��]�b]t�F���'-����������'-��x   x   F����q�b�X�P>�=�#���
�����	þ<��������z���g��a���g�#�z�����5����	þ~�边�
�>�#�P>�^�X��q�F����؋���쒿���؋�x   x   �q���Ki��9O��X4��5�(�D�ھ'k��������=�z���m���m�E�z�������2k��A�ھ(��5��X4��9O��Ki��q��'-����1���6�����$-��x   x   nu�L\���A���'� ��1��s˾,���{���.���{���u�!�{��.�����'����s˾+������'���A�L\�pu��L������쒿6���쒿�����L��x   x   y�d���K���1����w�دܾ~��Vj��������v~��v~������Hj��~��ܾ߯v������1���K�w�d�[7{���������������������\7{�x   x   ^�P��]8��> ���	�����`ɾ����e[��Z7����5���[7��p[�������`ɾ����	��> ��]8�g�P�Ccg�W7{��L��'-���؋�$-���L��\7{�Hcg�x   x   }j�q�m`�`�ξ�&��`5��Rz��O���ݭ�����᭍�M���Kz��[5���&��o�ξn`�p�tj�$���3�`�A��L��jS�~�U��jS��L�\�A���3�$�x   x   q�����Ҿ3I��gޭ��<��=:��,w��穏�婏�1w��@:���<��jޭ�I���Ҿ���u�!���> ���-���8�ީ@���D���D�ک@���8���-��> ���x   x   m`��Ҿ�
���а��椾,��[J��I钾?ϑ�H钾WJ��,���椾�а��
���Ҿf`�U? ���������#���+� M1�x!3��L1���+���#�������Z? �x   x   `�ξ3I���а��(���=���yS��U���^���zS����=���(���а�I��k�ξ@5��x��7���C����2��4����>�� ��2��x��35�x   x   �&��gޭ��椾�=��������������s��������������=���椾qޭ��&���ƾA�վ��0���(�R���x�����x�Q��(�=����B�վ%�ƾx   x   `5���<��,��������m���ꔾ�ꔾ�m�������,���<��\5�����挻��@Ǿ�\Ӿ��޾~�辜�������辺�޾�\Ӿ�@Ǿ،�����x   x   Rz��=:��[J��yS�������ꔾ픾�ꔾ����{S��fJ��;:��Lz��^@��i�������P��J���Rbƾ��̾ �о;	Ҿ/�о��̾SbƾW����P�����^���Z@��x   x   O���,w��I钾U����s���ꔾ�ꔾ�s��V���K钾(w��O������i����V������%%��N��d߭�(K��������'K��d߭�N��%�������V��t������x   x   ݭ��穏�?ϑ�^��������m������V���Bϑ�詏�ޭ��^7��O���P㋾�+��$A��"���1O������1������,������8O��$���,A���+��B㋾Q���_7��x   x   ���婏�H钾zS����������{S��K钾詏�����^�����׀������9��J�� ��)����:������ȕ���:������ ���I�2������ـ������^��x   x   ᭍�1w��WJ�������fJ��(w��ޭ���^�������{�	�r��wk���e���a�W_���]��(]��\��(]���]�W_���a���e��wk���r��{������^��x   x   M���@:��,���=���=��,��;:��O���^7������{���m�
�a�I�V��N��eG���B���?��'>��'>���?���B��eG��N�7�V��a���m�!�{����[7��x   x   Kz���<���椾�(���椾�<��Lz�����O���׀��	�r�
�a���Q��CD��'9�ș0���*�*'���%�,'���*�ߙ0��'9��CD���Q���a���r�΀��N������x   x   [5��jޭ��а��а�qޭ�\5��^@��i���P㋾�����wk�I�V��CD�{m4��'�����%p�p�������'�ym4��CD�>�V��wk�����G㋾h���e@��x   x   �&��I���
��I���&�����i����V���+��9����e��N��'9��'�������{�	� �s�	��������'��'9��N���e�(���+���V��e������x   x   o�ξ�Ҿ�Ҿk�ξ�ƾ挻��������$A��J���a��eG�ș0������f�>��I��T�}����Ι0�
fG���a�J�$A���������茻��ƾx   x   n`����f`�@5�A�վ�@Ǿ�P��%%��"���� ��W_���B���*���{�	�>��F��?��s�	�����*���B�W_�� ��(���%���P���@ǾF�վ;5�x   x   p�u�U? ��x�����\ӾJ���N��1O��)�����]���?�*'�%p� �I��?��# �p�'���?���]�%���6O��N��R����\Ӿ��y��W? �x   x   tj�!�����7�0�����޾Rbƾd߭������:���(]��'>���%�p�s�	�T�s�	�p���%��'>��(]��:������d߭�Rbƾ��޾0���7����!��x   x   $��> ������(�~�辢�̾)K��1�������\��'>�,'������}����'��'>��\�Ǖ��=�� K����̾x��(�!������> �$�x   x   ��3���-���#�C��R���� �о�������ȕ���(]���?���*����������*���?��(]�Ǖ���������,�о��P��>����#���-���3�6�x   x   `�A���8���+����x����;	Ҿ���,���:����]���B�ߙ0���'��'�Ι0���B���]��:��=�����<	Ҿ���x������+���8�^�A�xF�xF�x   x   �L�ީ@� M1�2��������/�о'K���������W_��eG��'9�ym4��'9�
fG�W_�%������� K��,�о��󾶹�0���L1�ݩ@�ݍL�wT�)�V�lT�x   x   �jS���D�x!3�4���x��𾔗̾d߭�8O��� ����a��N��CD��CD��N���a�� ��6O��d߭���̾��x�0��t!3���D��jS���]��:c��:c���]�x   x   ~�U���D��L1���Q�����SbƾN��$����I���e�7�V���Q�>�V���e�J�(���N��Rbƾx��P������L1���D�x�U���b�P3k�on�B3k���b�x   x   �jS�ک@���+�>��(���޾W���%��,A��2���wk��a���a��wk�'��$A��%��R�����޾(�>����+�ݩ@��jS���b���m���s�ʭs���m���b�x   x   �L���8���#� ��=����\Ӿ�P�������+��������r���m���r������+�������P���\Ӿ0���!����#���8�ݍL���]�P3k���s�F�v���s�H3k���]�x   x   \�A���-����2���@Ǿ����V��B㋾ـ���{�!�{�΀��G㋾�V������@Ǿ��7������-�^�A�wT��:c�on�ʭs���s�rn��:c�tT�x   x   ��3��> �����x��B�վ،��^���t���Q�������������N���h���e���茻�F�վy������> ���3�xF�)�V��:c�B3k���m�H3k��:c�!�V�xF�x   x   $���Z? �35�%�ƾ���Z@�����_7���^���^��[7�����e@������ƾ;5�W? �!��$�6�xF�lT���]���b���b���]�tT�xF�6�x   x   �$�#�۾�Wʾ�绾R���f5���l���מ��$���$���מ��l��[5��a����绾�Wʾ%�۾�$�p��R�#����!�%�'�H++�E++�%�'���!�#���R�r�x   x   #�۾-V̾s��uX��iޭ�$���lj��Ϡ��V��Ǡ��jj��0���jޭ�fX��s��3V̾%�۾���W? ��	���f��l��n4�l��d������	�V? ����x   x   �Wʾs�������а�̮��&���è�
,��	,���è�&��Ǯ���а�����s���Wʾ	q׾�#�y��v�PU�����N��N����OU�u�y���#�q׾x   x   �绾uX���а��������Z��N﫾'�N﫾^����������а�hX���绾8�ľ��ξ�^ھ��+��gw�����څ ����hw��&���}^ھ��ξ4�ľx   x   R���iޭ�̮������5��S g��g��P5������®��qޭ�`���'���D����¾%˾�\ӾA�ھ�߾�������߾:�ھ�\Ӿ%˾��¾�D��5��x   x   f5��$���&��Z��ScD��g���oD��MO��&��*���\5��`
��)t��[@��������R����	þ��žQ�ƾ��ž�	þM���������`@��t��f
��x   x   �l��lj���è�N﫾 g��g���d���g��V﫾�è�aj���l��^@���G�������?������@���N��|��������%|���M��F���ǯ���?�������G��T@��x   x   �מ�Ϡ��
,��'�g��oD��g��'�	,��Ơ���מ�r[��i������x����v|���W��6O������Q�����BO���W��r|�����x����o���f[��x   x   �$��V��	,��N﫾PMV﫾	,��T���$��T�����P㋾巇��������c��Ӏ�%���n���l���-���Ӏ��b���������𷇾B㋾��Y���x   x   �$��Ǡ���è�^��5��O���è�Ơ���$�������\���.�������v�(�m�w"g��|b�q�_���]��[]���]���_��|b��"g��m��v������.���\������x   x   �מ�jj��&����������&��aj���מ�T����\��%���B�z��wk�oe^�ܨS�OVK��UE�|A���?���?��{A��UE�KVK��S�}e^��wk�A�z�����\��R���x   x   �l��0���Ǯ�����®��*����l��r[�����.��B�z���g�I�V��H��<���2�M/,�O(�'�O(�?/,���2��<��H�L�V���g�E�z��.����p[��x   x   [5��jޭ��а��а�qޭ�\5��^@��i���P㋾�����wk�I�V��CD�{m4��'�����%p�p�������'�ym4��CD�>�V��wk�����G㋾h���e@��x   x   a���fX������hX��`���`
���G����巇��v�oe^��H�{m4�w�#������ ��!�# ������h�#�fm4��H�ve^���v���򓾐G��b
��x   x   �绾s��s���绾'��)t�������x�����(�m�ܨS��<��'�����D
�I��w�����?���D
�����'��<�ۨS��m�����x������&t��"��x   x   �Wʾ3V̾�Wʾ8�ľ�D��[@���?��������x"g�OVK���2�����I��&H����>H��I�������2�MVK�x"g��������?��`@���D��2�ľx   x   %�۾%�۾	q׾��ξ��¾�������v|��c���|b��UE�M/,��� �w����ڄ��� ����N/,��UE� }b��b��q|��ɯ�������¾��ξq׾x   x   �$𾝗�#澆^ھ%˾���@����W��Ӏ�q�_�|A�O(�%p��!����>H������!�%p�O(�|A�q�_�Ӏ��W��@������%˾�^ھ�#澝��x   x   p�W? �y�����\ӾR���N��6O��%�����]���?�'�p�# �?��I�� �%p�*'���?���]�)���1O��N��J����\Ӿ���x��U? �u�x   x   �R��	�v�+��A�ھ�	þ|�����n����[]���?�O(������D
������O(���?��[]�m������!|���	þD�ھ!��x���	��R����x   x   #����PU�gw���߾��ž����Q��l�����]��{A�?/,�����������N/,�|A���]�m����Q�������ž�߾ow��MU���"���Q��Q�x   x   ��!�f�����������Q�ƾ������-�����_��UE���2���'�h�#��'��2��UE�q�_�)���������B�ƾ��⾃�����i��}�!��;'�/0)��;'�x   x   %�'�l���N�څ ������ž%|��BO��Ӏ��|b�KVK��<�ym4�fm4��<�MVK� }b�Ӏ�1O��!|����ž���ۅ ��N�i��'�'�0�/�:�3�;�3�0�/�x   x   H++�n4��N�����߾�	þ�M���W���b���"g��S��H��CD��H�ۨS�x"g��b���W��N���	þ�߾����N�u4�C++�h95�h�;��=�o�;�g95�x   x   E++�l�����hw��:�ھM���F���r|�������m�}e^�L�V�>�V�ve^��m�����q|��@���J���D�ھow�����i��C++�K7�O�?�*D�(D�M�?�M7�x   x   %�'�d��OU�&���\Ӿ���ǯ��������v��wk���g��wk���v������ɯ������\Ӿ!��MU�i��'�'�h95�O�?��2F��tH��2F�S�?�h95�x   x   ��!���u��%˾����?���x��𷇾����A�z�E�z�������x���?�����%˾��x���}�!�0�/�h�;�*D��tH��tH�(D�h�;�1�/�x   x   #����	�y��}^ھ��¾`@��������B㋾�.������.��G㋾�򓾯���`@����¾�^ھ�x����	�"���;'�:�3��=�(D��2F�(D�#�=�9�3��;'�x   x   �R�V? ��#澇�ξ�D��t���G��o������\���\����h����G��&t���D����ξ�#�U? ��R��Q�/0)�;�3�o�;�M�?�S�?�h�;�9�3�10)��Q�x   x   r����q׾4�ľ5��f
��T@��f[��Y�������R���p[��e@��b
��"��2�ľq׾���u�����Q��;'�0�/�g95�M7�h95�1�/��;'��Q����x   x   7�о�Ǿ�����绾�&��@ط��o��|l��(v��l���o��6ط��&���绾�����Ǿ1�о%�۾n`辣$���u �O5�J�h[	�J�R5��u ��$��q`�&�۾x   x   �Ǿ={¾s��1I��yr��?R���O��u���u����O��GR���r��I��s��C{¾�Ǿ`�ξq׾;5���꾒�����Bb��Vb������������<5�q׾Y�ξx   x   ����s���
��I���3Wľ�ƾQjȾ�ɾMjȾ�ƾ&WľJ����
��s��������þȾ��ξF�վܾ߯�_⾤&�Oy羝&澒_��ܾB�վ��ξɏȾ��þx   x   �绾1I��I���>ƾʾ7;��ξ��ξ7;ʾHƾC���I���绾T4��	=���ﾾ��¾�@Ǿ�s˾��ξ�о�о��ξ�s˾�@Ǿ��¾�ﾾ=��N4��x   x   �&��yr��3Wľʾ��ξ�Ҿ;.Ӿ�Ҿ��ξʾ+Wľ�r���&��'�������±��j������P��2k��빾�u��빾$k���P������j���±�����,��x   x   @ط�?R���ƾ7;�Ҿ��Ծ��Ծ�Ҿ
7;�ƾJR��:ط����)t���\��褾�̣�ɯ��%��5����$���$��;���%%��Ư���̣�	褾�\��t�����x   x   �o���O��QjȾ��ξ;.Ӿ��Ծ?.Ӿ��ξNjȾ�O���o������i��������H��np����q|��(����s���`���s��#���k|����wp���H������]�������x   x   |l��u����ɾ��ξ�Ҿ�Ҿ��ξ�ɾt����l��R��Jj���V���x�����9��\����b��� ���~�0�~�� ���b��b����8������x���V��[j��R��x   x   (v��v���MjȾ7;��ξ
7;NjȾt���$v���Ȭ�,�������+������,{��p�+�g� }b�W_�qQ^�W_��|b�$�g��p��,{�����+����.����Ȭ�x   x   l���O���ƾʾʾ�ƾ�O���l���Ȭ��0���l�����9��(�m�7�^��RS���J��UE���B���B��UE���J��RS�/�^��m�2������l���0���Ȭ�x   x   �o��GR��&WľHƾ+WľJR���o��R��,����l�� ���z���e�ܨS���D�<,9�`1�N/,���*�[/,�M1�B,9���D��S���e��z����l��(���R��x   x   6ط��r��J���C����r��:ط�����Jj���������z�<@c��N��<��t-���"�Q>������j>���"��t-��<�~N�=@c�#�z�������Hj������x   x   �&��I���
��I���&�����i����V���+��9����e��N��'9��'�������{�	� �s�	��������'��'9��N���e�(���+���V��e������x   x   �绾s��s���绾'��)t�������x�����(�m�ܨS��<��'�����D
�I��w�����?���D
�����'��<�ۨS��m�����x������&t��"��x   x   ����C{¾����T4�������\���H������,{�7�^���D��t-�����D
�������ڄ�F���D
���� u-���D�6�^��,{�����H���\������U4��x   x   �Ǿ�Ǿ��þ	=���±�褾np��9���p��RS�<,9���"����I������r����>�������"�8,9��RS��p��8��rp��	褾�±�=����þx   x   1�о`�ξȾ�ﾾ�j���̣���\���+�g���J�`1�Q>�{�	�w�����r�潵��w��{�	�Q>�`1���J�+�g�\������̣��j���ﾾȾ`�ξx   x   %�۾q׾��ξ��¾���ɯ��q|���b�� }b��UE�N/,���� ����ڄ���w�� ���M/,��UE��|b�c��v|�����������¾��ξ	q׾%�۾x   x   n`�;5�F�վ�@Ǿ�P��%��(���� ��W_���B���*���s�	�?��F��>��{�	�����*���B�W_�� ��"���%%���P���@ǾA�վ@5�f`����x   x   �$�����ܾ߯�s˾2k��5����s���~�qQ^���B�[/,�j>�����D
��D
����Q>�M/,���B�|Q^�$�~��s��/���)k���s˾�ܾ��꾣$��w��w��x   x   �u ����_⾥�ξ빾�$���`��0�~�W_��UE�N1���"������������"�`1��UE�W_�$�~��`���$��)빾��ξ�_⾎���u �H��d+�A��x   x   O5������&��о�u���$���s��� ���|b���J�B,9��t-��'��'� u-�8,9���J��|b�� ���s���$���u���о�&澍���U5���I.�N.���x   x   J�Bb��Oy��о빾;���#����b��$�g��RS���D��<��'9��<���D��RS�+�g�c��"���/���)빾�оUy�Jb��J������$�����x   x   h[	�Vb���&澪�ξ$k��%%��k|��b����p�/�^��S�}N��N�ۨS�6�^��p�\���v|��%%��)k����ξ�&�Jb��h[	�9�v��U��U��v��9�x   x   J������_⾐s˾�P��Ư�����8���,{��m���e�=@c���e��m��,{��8���𓾹����P���s˾�_⾍���J�9�Y������� ����Z��9�x   x   R5�����ܾ�@Ǿ����̣�wp��������2���z�#�z�'��������rp���̣�����@Ǿ�ܾ���U5���v�����z6"�w6"����z����x   x   �u ����B�վ��¾�j��	褾�H���x���+�����������+���x���H��	褾�j����¾A�վ����u �����U���� �w6"��� �Q������x   x   �$��<5ᾈ�ξ�ﾾ�±��\�������V�����l���l������V�������\���±��ﾾ��ξ@5ᾣ$��H��I.��$�U��������Q���$�L.�F��x   x   q`�q׾ɏȾ=������t��]���[j��.����0��(���Hj��e���&t������=��Ⱦ	q׾f`�w��d+�N.���v��Z��z����L.�c+�w��x   x   &�۾Y�ξ��þN4��,���������R���Ȭ��Ȭ�R���������"��U4����þ`�ξ%�۾���w��A������9�9�����F��w�����x   x   g�ƾ�Ǿ�Wʾf�ξ@`Ӿ2�׾��۾��ݾ��ݾ��۾(�׾X`Ӿo�ξ�Wʾ�Ǿ\�ƾ�Ǿ�Wʾo�ξX`Ӿ(�׾��۾��ݾ��ݾ��۾2�׾@`Ӿf�ξ�Wʾ�Ǿx   x   �Ǿ(V̾�Ҿ��پH���c��<�����<��c�F�ྗ�پ�Ҿ3V̾�ǾȠľ��þ2�ľ�ƾ�`ɾ�˾�;x�ξ#�;��˾�`ɾ$�ƾ3�ľ��þ��ľx   x   �Wʾ�Ҿ;�۾?徢C�&Z�ݙ��ԙ��Z�C�E�J�۾�Ҿ�Wʾ��þ=���=���D��茻�~��у��'��'��΃��~��ڌ���D��=��A�����þx   x   f�ξ��پ?�{��r ��,������=���l ��x��<從�پk�ξ8�ľ	=�������±�`@�����'�������옭�����-������a@��ñ�����=��3�ľx   x   @`ӾH�ྡྷC�r ���	 ��"��"�|	 �} ���C�I��Q`Ӿ�ƾ�D���±��M��	褾�?���������-��-��
��������?���社�M��ñ��D��$�ƾx   x   2�׾�c�&Z�,����"��F��"�1���Z��c�)�׾�`ɾ挻�[@��褾����rp����$A�������-������.A����sp�������社a@��ڌ���`ɾx   x   ��۾�<�ݙ������"��"����љ���<꾞�۾��˾~������?��np��vȍ��8������J��u|��u|�J������8��|ȍ�sp���?�����~����˾x   x   ��ݾ���ԙ��=���|	 �1���љ���뾤�ݾ#�;Ӄ�����������9��,$}��p�x"g���a��*`���a�w"g��p�*$}��8��������-���΃��#�;x   x   ��ݾ�<�Z�l ��} ��Z��<꾤�ݾy�ξ'���������$A�������p�{�_��RS�MVK�
fG��eG�MVK��RS�i�_��p�����.A��
�������'��x�ξx   x   ��۾�c澪C�x�ﾞC��c澞�۾#�;'��ۘ��-������J�w"g��RS��D�8,9��2�Ι0���2�B,9��D��RS�w"g�J�����-��옭�'���;x   x   (�׾F��E�<�I��)�׾��˾Ӄ������-���-��yu|���a�OVK�<,9���+���"�������"�}�+�B,9�MVK���a��u|��-��-������у���˾x   x   X`Ӿ��پJ�۾��پQ`Ӿ�`ɾ~������������yu|��*`��eG���2���"���������}�������"���2��eG��*`��u|��������'���~���`ɾx   x   o�ξ�Ҿ�Ҿk�ξ�ƾ挻��������$A��J���a��eG�ș0������f�>��I��T�}����Ι0�
fG���a�J�$A���������茻��ƾx   x   �Wʾ3V̾�Wʾ8�ľ�D��[@���?��������w"g�OVK���2�����I��&H����>H��I�������2�MVK�x"g��������?��`@���D��2�ľx   x   �Ǿ�Ǿ��þ	=���±�褾np��9���p��RS�<,9���"����I������r����>�������"�8,9��RS��p��8��rp��	褾�±�=����þx   x   \�ƾȠľ=��������M������vȍ�,$}�{�_��D���+����f�&H�����).⽓��&H��f������+��D�{�_�,$}�vȍ������M������=���Ƞľx   x   �Ǿ��þ=���±�	褾rp���8���p��RS�9,9���"����>����r�潓����I�������"�<,9��RS��p�9��np��褾�±�	=����þ�Ǿx   x   �Wʾ2�ľ�D��`@���?��������x"g�MVK��2�����I��>H����&H��I��������2�OVK�w"g��������?��[@���D��8�ľ�Wʾ3V̾x   x   o�ξ�ƾ茻��������$A��J���a�
fG�Ι0���}��T�I��>��f������ș0��eG���a�J�$A���������挻��ƾk�ξ�Ҿ�Ҿx   x   X`Ӿ�`ɾ~��'�����������u|��*`��eG���2���"����}������������"���2��eG��*`�yu|�����������~���`ɾQ`Ӿ��پJ�۾��پx   x   (�׾�˾у������-���-���u|���a�MVK�B,9�}�+���"�������"���+�<,9�OVK���a�yu|��-��-������Ӄ����˾)�׾I��<�E�F��x   x   ��۾�;'��옭�-������J�w"g��RS��D�B,9���2�Ι0��2�8,9��D��RS�w"g�J�����-��ۘ��'��#�;��۾�c澞C�x�ﾪC��c�x   x   ��ݾx�ξ'������
���.A�������p�i�_��RS�MVK��eG�
fG�MVK��RS�{�_��p�����$A���������'��y�ξ��ݾ�<�Z�} ��l ��Z��<�x   x   ��ݾ#�;΃��-����������8��*$}��p�w"g���a��*`���a�x"g��p�,$}�9�����������Ӄ��#�;��ݾ��љ��1���|	 �=���ԙ�����x   x   ��۾��˾~������?��sp��|ȍ��8������J��u|��u|�J������8��vȍ�np���?�����~����˾��۾�<�љ������"��"����ݙ���<�x   x   2�׾�`ɾڌ��a@���社����sp����.A�������-������$A����rp������褾Z@��挻��`ɾ)�׾�c�Z�1����"��F��"�,���&Z��c�x   x   @`Ӿ$�ƾ�D��ñ��M���社�?������
���-��-����������?��	褾�M���±��D���ƾQ`ӾI�ྞC�} ��|	 ��"��"��	 �r ���C�H��x   x   f�ξ3�ľ=������ñ�a@�����-�������옭�����'������`@���±�����	=��8�ľk�ξ��پ<�x��l ��=������,���r ��{��?循�پx   x   �Wʾ��þA���=���D��ڌ��~��΃��'��'��у��~��茻��D��=��=�����þ�Wʾ�ҾJ�۾E循C�Z�ԙ��ݙ��&Z�C�?�;�۾�Ҿx   x   �Ǿ��ľ��þ3�ľ$�ƾ�`ɾ��˾#�;x�ξ�;�˾�`ɾ�ƾ2�ľ��þȠľ�Ǿ3V̾�Ҿ��پF���c��<�����<��c�H�ྪ�پ�Ҿ(V̾x   x   7�о&�۾q`辠$���u �R5�J�h[	�J�O5��u ��$��n`�%�۾1�о�Ǿ�����绾�&��6ط��o��l��(v��|l���o��@ط��&���绾�����Ǿx   x   &�۾���w��F������9�9�����A��w�����%�۾`�ξ��þU4��"���������R���Ȭ��Ȭ�R���������,��N4����þY�ξx   x   q`�w��b+�L.���z��Z��v����N.�d+�w��f`�	q׾Ⱦ=������&t��e���Hj��(����0��.���[j��]���t������=��ɏȾq׾x   x   �$��F��L.��$�Q��������U���$�I.�H���$��@5ᾊ�ξ�ﾾ�±��\�������V������l���l�����V�������\���±��ﾾ��ξ<5�x   x   �u �����Q���� �w6"��� �U�������u ����A�վ��¾�j��	褾�H���x���+�����������+���x���H��	褾�j����¾B�վ���x   x   R5���z�����w6"�z6"����v����U5�����ܾ�@Ǿ����̣�rp��������(��#�z��z�2��������wp���̣�����@Ǿ�ܾ���x   x   J�9�Z������� ����Y��9�J������_⾇s˾�P���������8���,{��m���e�=@c���e��m��,{��8����Ư���P���s˾�_⾐���x   x   h[	�9�v��U��U��v��9�h[	�Jb���&澤�ξ)k��%%��v|��\����p�6�^�ۨS��N�}N��S�/�^��p�b���k|��%%��$k����ξ�&�Vb��x   x   J������$�����J�Jb��Uy��о)빾/���"���c��+�g��RS���D��<��'9��<���D��RS�$�g��b��#���;���빾�оOy�Bb��x   x   O5���N.�I.���U5������&��о�u���$���s��� ���|b���J�8,9� u-��'��'��t-�B,9���J��|b�� ���s���$���u���о�&澉���x   x   �u �A��d+�H���u ����_⾤�ξ)빾�$���`��$�~�W_��UE�`1���"������������"�M1��UE�W_�0�~��`���$��빾��ξ�_⾒��x   x   �$��w��w���$������ܾ�s˾)k��/����s��$�~�|Q^���B�M/,�Q>�����D
��D
����j>�[/,���B�qQ^��~��s��5���2k���s˾ܾ߯���x   x   n`����f`�@5�A�վ�@Ǿ�P��%%��"���� ��W_���B���*���{�	�>��F��?��s�	�����*���B�W_�� ��(���%���P���@ǾF�վ;5�x   x   %�۾%�۾	q׾��ξ��¾�������v|��c���|b��UE�M/,��� �w����ڄ��� ����N/,��UE� }b��b��q|��ɯ�������¾��ξq׾x   x   1�о`�ξȾ�ﾾ�j���̣���\���+�g���J�`1�Q>�{�	�w�����r�潵��w��{�	�Q>�`1���J�+�g�\������̣��j���ﾾȾ`�ξx   x   �Ǿ��þ=���±�	褾rp���8���p��RS�9,9���"����>����r�潓����I�������"�<,9��RS��p�9��np��褾�±�	=����þ�Ǿx   x   ����U4�������\���H������,{�6�^���D� u-�����D
�F��ڄ��������D
�����t-���D�7�^��,{�����H���\������T4������C{¾x   x   �绾"��&t�������x������m�ۨS��<��'�����D
�?�����w��I���D
�����'��<�ܨS�(�m�����x������)t��'���绾s��s��x   x   �&�����e����V���+��(����e��N��'9��'�������s�	� �{�	��������'��'9��N���e�9���+���V��i�������&��I���
��I��x   x   6ط�����Hj��������#�z�=@c�~N��<��t-���"�j>������Q>���"��t-��<��N�<@c��z�������Jj������:ط��r��C���J����r��x   x   �o��R��(����l�����z���e��S���D�B,9�M1�[/,���*�N/,�`1�<,9���D�ܨS���e��z� ���l��,���R���o��JR��+WľHƾ&WľGR��x   x   l���Ȭ��0���l�����2���m�/�^��RS���J��UE���B���B��UE���J��RS�7�^�(�m�9������l���0���Ȭ��l���O���ƾʾʾ�ƾ�O��x   x   (v���Ȭ�.������+������,{��p�$�g��|b�W_�qQ^�W_� }b�+�g��p��,{�����+�����,����Ȭ�$v��t���NjȾ
7;��ξ7;MjȾv���x   x   |l��R��[j���V���x������8��b����b��� ��0�~��~�� ���b��\���9������x���V��Jj��R���l��t����ɾ��ξ�Ҿ�Ҿ��ξ�ɾu���x   x   �o������]��������H��wp����k|��#����s���`���s��(���q|����np���H������i��������o���O��NjȾ��ξ?.Ӿ��Ծ;.Ӿ��ξQjȾ�O��x   x   @ط����t���\��	褾�̣�Ư��%%��;����$���$��5���%��ɯ���̣�褾�\��)t�����:ط�JR���ƾ
7;�Ҿ��Ծ��Ծ�Ҿ7;�ƾ?R��x   x   �&��,�������±��j������P��$k��빾�u��빾2k���P������j���±�����'���&���r��+Wľʾ��ξ�Ҿ;.Ӿ�Ҿ��ξʾ3Wľyr��x   x   �绾N4��=���ﾾ��¾�@Ǿ�s˾��ξ�о�о��ξ�s˾�@Ǿ��¾�ﾾ	=��T4���绾I��C���Hƾʾ7;��ξ��ξ7;ʾ>ƾI���1I��x   x   ������þɏȾ��ξB�վ�ܾ�_⾝&�Oy群&澐_�ܾ߯F�վ��ξȾ��þ����s���
��J���&Wľ�ƾMjȾ�ɾQjȾ�ƾ3WľI����
��s��x   x   �ǾY�ξq׾<5���꾑�����Vb��Bb������������;5�q׾`�ξ�ǾC{¾s��I���r��GR���O��u���u����O��?R��yr��1I��s��={¾x   x   �$�r��R�#����!�%�'�E++�H++�%�'���!�#���R�p��$�%�۾�Wʾ�绾a���[5���l���מ��$���$���מ��l��f5��R����绾�Wʾ#�۾x   x   r�����Q��;'�1�/�h95�M7�g95�0�/��;'��Q����u����q׾2�ľ"��b
��e@��p[��R�������Y���f[��T@��f
��5��4�ľq׾���x   x   �R��Q�10)�9�3�h�;�S�?�M�?�o�;�;�3�/0)��Q��R�U? ��#澐�ξ�D��&t���G��h������\���\����o����G��t���D����ξ�#�V? �x   x   #���;'�9�3�#�=�(D��2F�(D��=�:�3��;'�"����	��x���^ھ��¾`@��������G㋾�.������.��B㋾�򓾴���`@����¾}^ھy����	�x   x   ��!�1�/�h�;�(D��tH��tH�*D�h�;�0�/�}�!���x���%˾����?���x�������E�z�A�z�����𷇾�x���?�����%˾�u���x   x   %�'�h95�S�?��2F��tH��2F�O�?�h95�'�'�i��MU�!���\Ӿ���ɯ���������v��wk���g��wk��v������ǯ������\Ӿ&��OU�d��x   x   E++�M7�M�?�(D�*D�O�?�L7�C++�i�����ow��D�ھJ���@���q|�������m�ve^�>�V�L�V�}e^��m�����r|��F���M���:�ھhw�����l��x   x   H++�g95�o�;��=�h�;�h95�C++�u4��N�����߾�	þN���W���b��x"g�ۨS��H��CD��H��S��"g��b���W���M���	þ�߾����N�n4�x   x   %�'�0�/�;�3�:�3�0�/�'�'�i���N�ۅ ������ž!|��1O��Ӏ� }b�MVK��<�fm4�ym4��<�KVK��|b�Ӏ�BO��%|����ž���څ ��N�l��x   x   ��!��;'�/0)��;'�}�!�i�����������B�ƾ������)���q�_��UE��2��'�h�#���'���2��UE���_�-���������Q�ƾ��⾅�����f��x   x   #���Q��Q�"����MU�ow���߾��ž����Q��m�����]�|A�N/,�����������?/,��{A���]�l����Q�������ž�߾gw��PU���x   x   �R�����R���	�x�!��D�ھ�	þ!|�����m����[]���?�O(�������D
�����O(���?��[]�n������|���	þA�ھ+��v��	�x   x   p�u�U? ��x�����\ӾJ���N��1O��)�����]���?�*'�%p� �I��?��# �p�'���?���]�%���6O��N��R����\Ӿ��y��W? �x   x   �$𾝗�#澆^ھ%˾���@����W��Ӏ�q�_�|A�O(�%p��!����>H������!�%p�O(�|A�q�_�Ӏ��W��@������%˾�^ھ�#澝��x   x   %�۾q׾��ξ��¾���ɯ��q|���b�� }b��UE�N/,���� ����ڄ���w�� ���M/,��UE��|b�c��v|�����������¾��ξ	q׾%�۾x   x   �Wʾ2�ľ�D��`@���?��������x"g�MVK��2�����I��>H����&H��I��������2�OVK�w"g��������?��[@���D��8�ľ�Wʾ3V̾x   x   �绾"��&t�������x������m�ۨS��<��'�����D
�?�����w��I���D
�����'��<�ܨS�(�m�����x������)t��'���绾s��s��x   x   a���b
���G�������v�ve^��H�fm4�h�#������# ��!� ������w�#�{m4��H�oe^��v�巇��򓾗G��`
��`���hX������fX��x   x   [5��e@��h���G㋾�����wk�>�V��CD�ym4���'�����p�%p������'�{m4��CD�I�V��wk�����P㋾i���^@��\5��qޭ��а��а�jޭ�x   x   �l��p[�����.��E�z���g�L�V��H��<���2�?/,�O(�'�O(�M/,���2��<��H�I�V���g�B�z��.����r[���l��*���®�����Ǯ��0���x   x   �מ�R����\�����A�z��wk�}e^��S�KVK��UE��{A���?���?�|A��UE�OVK�ܨS�oe^��wk�B�z�$����\��T����מ�aj��&����������&��jj��x   x   �$�������\���.�������v��m��"g��|b���_���]��[]���]�q�_��|b�w"g�(�m��v������.���\�������$��Ơ���è�O��5��^���è�Ǡ��x   x   �$��Y�����B㋾𷇾��������b��Ӏ�-���l���n���%���Ӏ�c���������巇�P㋾��T����$��T��	,��V﫾MPN﫾	,��V��x   x   �מ�f[��o������x����r|���W��BO������Q�����6O���W��v|�����x����i���r[���מ�Ơ��	,��'�g��oD��g��'�
,��Ϡ��x   x   �l��T@���G�������?��ǯ��F����M��%|��������|��N��@��������?�������G��^@���l��aj���è�V﫾g��d���g��� g��N﫾�è�lj��x   x   f5��f
��t��`@��������M����	þ��žQ�ƾ��ž�	þR���������Z@��)t��`
��\5��*���&��O��MoD��g���cD��SZ��&��$���x   x   R���5���D����¾%˾�\Ӿ:�ھ�߾�������߾A�ھ�\Ӿ%˾��¾�D��'��`���qޭ�®������5��Pg�� g��S5������̮��iޭ�x   x   �绾4�ľ��ξ}^ھ�&��hw�����څ ����gw��+���澆^ھ��ξ8�ľ�绾hX���а��������^��N﫾'�N﫾Z����������а�uX��x   x   �Wʾq׾�#�y��u�OU�����N��N����PU�v�y���#�	q׾�Wʾs�������а�Ǯ��&���è�	,��
,���è�&��̮���а�����s��x   x   #�۾���V? ���	���d��l��n4�l��f�����	�W? ����%�۾3V̾s��fX��jޭ�0���jj��Ǡ��V��Ϡ��lj��$���iޭ�uX��s��-V̾x   x   }j�$���3�\�A��L��jS�~�U��jS��L�`�A���3�$�tj�p�n`�o�ξ�&��[5��Kz��M���᭍����ݭ��O���Rz��`5���&��`�ξm`�q�x   x   $�6�xF�tT���]���b���b���]�lT�xF�6�$�!��W? �;5��ƾ���e@�����[7���^���^��_7�����Z@�����%�ƾ35�Z? ���x   x   ��3�xF�!�V��:c�H3k���m�B3k��:c�)�V�xF���3��> ����y��F�վ茻�e���h���N�������������Q���t���^���،��B�վ�x������> �x   x   \�A�tT��:c�rn���s�ʭs�on��:c�wT�^�A���-����7����@Ǿ����V��G㋾΀��!�{��{�ـ��B㋾�V������@Ǿ�2������-�x   x   �L���]�H3k���s�F�v���s�P3k���]�ݍL���8���#�!��0����\Ӿ�P�������+��������r���m���r������+�������P���\Ӿ=��� ����#���8�x   x   �jS���b���m�ʭs���s���m���b��jS�ݩ@���+�>��(���޾R���%��$A��'���wk���a��a��wk�2��,A��%��W�����޾(�>����+�ک@�x   x   ~�U���b�B3k�on�P3k���b�x�U���D��L1����P��x��RbƾN��(���J���e�>�V���Q�7�V���e��I�$���N��Sbƾ���Q�����L1���D�x   x   �jS���]��:c��:c���]��jS���D�t!3�0��x��𾤗̾d߭�6O��� ����a��N��CD��CD��N���a�� ��8O��d߭���̾��x�4��x!3���D�x   x   �L�lT�)�V�wT�ݍL�ݩ@��L1�0��������,�о K������%���W_�
fG��'9�ym4��'9��eG�W_��������'K��/�о��󾰹�2�� M1�ީ@�x   x   `�A�xF�xF�^�A���8���+����x����<	Ҿ���=���:����]���B�Ι0��'���'�ߙ0���B���]��:��,�����;	Ҿ���x�����+���8�x   x   ��3�6���3���-���#�>��P����,�о�������Ǖ���(]���?���*����������*���?��(]�ȕ��������� �о��R��C����#���-�x   x   $�$��> ����!��(�x�辤�̾ K��=��Ǖ���\��'>�'���}�������,'��'>��\�����1��(K����̾~��(�������> �x   x   tj�!�����7�0�����޾Rbƾd߭������:���(]��'>���%�p�s�	�T�s�	�p���%��'>��(]��:������d߭�Rbƾ��޾0���7����!��x   x   p�W? �y�����\ӾR���N��6O��%�����]���?�'�p�# �?��I�� �%p�*'���?���]�)���1O��N��J����\Ӿ���x��U? �u�x   x   n`�;5�F�վ�@Ǿ�P��%��(���� ��W_���B���*���s�	�?��F��>��{�	�����*���B�W_�� ��"���%%���P���@ǾA�վ@5�f`����x   x   o�ξ�ƾ茻��������$A��J���a�
fG�Ι0���}��T�I��>��f������ș0��eG���a�J�$A���������挻��ƾk�ξ�Ҿ�Ҿx   x   �&�����e����V���+��(����e��N��'9��'�������s�	� �{�	��������'��'9��N���e�9���+���V��i�������&��I���
��I��x   x   [5��e@��h���G㋾�����wk�>�V��CD�ym4���'�����p�%p������'�{m4��CD�I�V��wk�����P㋾i���^@��\5��qޭ��а��а�jޭ�x   x   Kz�����N���΀����r���a���Q��CD��'9�ߙ0���*�,'���%�*'���*�ș0��'9��CD���Q�
�a�	�r�׀��O������Lz���<���椾�(���椾�<��x   x   M���[7�����!�{���m��a�7�V��N��eG���B���?��'>��'>���?���B��eG��N�I�V�
�a���m��{����^7��O���;:��,���=���=��,��@:��x   x   ᭍��^�������{���r��wk���e���a�W_���]��(]��\��(]���]�W_���a���e��wk�	�r��{������^��ޭ��(w��fJ�������WJ��1w��x   x   ����^�����ـ������2���I�� ������:��ȕ�������:��)���� ��J�9������׀������^�����詏�K钾{S����������zS��H钾婏�x   x   ݭ��_7��Q���B㋾�+��,A��$���8O������,������1������1O��"���$A���+��P㋾O���^7��ޭ��詏�Bϑ�V��������m������^���?ϑ�穏�x   x   O������t����V������%��N��d߭�'K��������(K��d߭�N��%%�������V��i������O���(w��K钾V����s���ꔾ�ꔾ�s��U���I钾,w��x   x   Rz��Z@��^�������P��W���Sbƾ��̾.�о;	Ҿ �о��̾RbƾJ����P�����i���^@��Lz��;:��fJ��{S�������ꔾ픾�ꔾ����yS��[J��=:��x   x   `5�����،���@Ǿ�\Ӿ��޾��辟������~����޾�\Ӿ�@Ǿ挻����\5���<��,��������m���ꔾ�ꔾ�m�������,���<��x   x   �&��%�ƾB�վ�=���(�Q���x�����x�R��(�0�����A�վ�ƾ�&��qޭ��椾�=��������������s��������������=���椾gޭ�x   x   `�ξ35��x��2� ��>����4��2����C����7��x��@5�k�ξI���а��(���=���zS��^���U���yS����=���(���а�3I��x   x   m`�Z? ���������#���+��L1�x!3� M1���+���#�������U? �f`��Ҿ�
���а��椾,��WJ��H钾?ϑ�I钾[J��,���椾�а��
���Ҿx   x   q����> ���-���8�ک@���D���D�ީ@���8���-��> �!��u�����ҾI��jޭ��<��@:��1w��婏�穏�,w��=:���<��gޭ�3I���Ҿ���x   x   O�:�^�P�y�d�nu��q��F���I����q��ju���d�_�P�G�:�$��R��$��X`Ӿ6ط��l��M���L���>���8���Q���J����l��Bط�F`Ӿ�$���R�$�x   x   ^�P�Hcg�\7{��L��$-���؋�'-���L��W7{�Ccg�g�P��]8��> ��	���꾼`ɾ����p[��[7����5���Z7��e[�������`ɾ�����	��> ��]8�x   x   y�d�\7{���������������������[7{�w�d���K���1����v�ܾ߯~��Hj��������v~��v~������Vj��~��دܾw������1���K�x   x   nu��L������쒿6���쒿�����L��pu�L\���A���'���+��s˾'�������.��!�{���u��{��.��{��,����s˾1�� ����'���A�L\�x   x   �q��$-����6���1�����'-���q���Ki��9O��X4��5�(�A�ھ2k��������E�z���m���m�=�z�������'k��D�ھ(��5��X4��9O��Ki�x   x   F����؋���쒿���؋�F����q�^�X�P>�>�#���
�~���	þ5�������#�z���g��a���g��z�����<����	þ��辷�
�=�#�P>�b�X��q�x   x   I���'-����������'-��F���b]t��]���D���*���������̾|���s���u|�=@c�L�V�7�V�N@c�}u|��s��|����̾��������*���D��]�d]t�x   x   �q���L�������L���q���q��]�{�F��c.��������%5Ծ(K������~��*`�}N��H��N��*`�2�~����+K��%5Ծ~�������c.�y�F��]��q�x   x   ju�W7{�[7{�pu��Ki�^�X���D��c.� i�v� پ���1��n���qQ^��eG��<��<��eG�`Q^�i���0�����( پw��h��c.���D�d�X��Ki�x   x   ��d�Ccg�w�d�L\��9O�P>���*����v���ھ�ַ����������[]���B���2��t-���2���B��[]�ƕ�������ַ�{�ھr������*�P>��9O�L\�x   x   _�P�g�P���K���A��X4�>�#������� پ�ַ������%���\���?�[/,���"���"�?/,���?�
�\��%�������ַ�# پ������=�#��X4���A���K�x   x   G�:��]8���1���'��5���
�����%5Ծ��������%����\��'>�O(�j>����j>�O(��'>���\��%���������%5Ծ������
��5���'���1��]8�x   x   $��> ������(�~�辢�̾(K��1�������\��'>�,'������}����'��'>��\�Ǖ��=�� K����̾x��(�!������> �$�x   x   �R��	�v�+��A�ھ�	þ|�����n����[]���?�O(������D
������O(���?��[]�m������!|���	þD�ھ!��x���	��R����x   x   �$�����ܾ߯�s˾2k��5����s���~�qQ^���B�[/,�j>�����D
��D
����Q>�M/,���B�|Q^�$�~��s��/���)k���s˾�ܾ��꾣$��w��w��x   x   X`Ӿ�`ɾ~��'�����������u|��*`��eG���2���"����}������������"���2��eG��*`�yu|�����������~���`ɾQ`Ӿ��پJ�۾��پx   x   6ط�����Hj��������#�z�=@c�~N��<��t-���"�j>������Q>���"��t-��<��N�<@c��z�������Jj������:ط��r��C���J����r��x   x   �l��p[�����.��E�z���g�L�V��H��<���2�?/,�O(�'�O(�M/,���2��<��H�I�V���g�B�z��.����r[���l��*���®�����Ǯ��0���x   x   M���[7�����!�{���m��a�7�V��N��eG���B���?��'>��'>���?���B��eG��N�I�V�
�a���m��{����^7��O���;:��,���=���=��,��@:��x   x   L�����v~���u���m���g�N@c��*`�`Q^��[]�
�\���\��\��[]�|Q^��*`�<@c���g���m���u��v~��K���jΌ�n-���[�����[��j-��fΌ�x   x   >����5���v~��{�=�z��z�}u|�2�~�i���ƕ���%���%��Ǖ��m���$�~�yu|��z�B�z��{��v~��5��:���X���j��.-��-!��.!��2-���j��W��x   x   8��������.����������s�����0��������������=������s����������.������:���.郾�����f��� ��2:��� ���f������0郾x   x   Q���Z7����{�����<���|��*K������ַ��ַ���� K��!|��/�����������^7��K���X������9Ճ�����h��h������4Ճ�����\��x   x   J���e[��Vj��,���'k���	þ��̾%5Ծ( پ{�ھ# پ%5Ծ��̾�	þ)k�����Jj��r[��O���jΌ��j���f�������|��o+���|�������f���j��eΌ�x   x   �l������~���s˾D�ھ�������~���w�r���������x��D�ھ�s˾~�������l��;:��n-��.-��� ��h��o+��r+��h��� ��2-��q-��<:��x   x   Bط��`ɾدܾ1��(���
�������h��������
�(�!���ܾ�`ɾ:ط�*���,���[��-!��2:��h���|��h��0:��/!���[��,��&���x   x   F`Ӿ���w� ���5�=�#���*��c.��c.���*�=�#��5�!��x����Q`Ӿ�r��®���=����.!��� ����������� ��/!�����=��̮��}r��x   x   �$����	������'��X4�P>���D�y�F���D�P>��X4���'������	��$����پC�������=���[��2-���f��4Ճ��f��2-���[���=�����H�����پx   x   �R��> ���1���A��9O�b�X��]��]�d�X��9O���A���1��> ��R�w��J�۾J���Ǯ��,��j-���j�����������j��q-��,��̮��H���2�۾w��x   x   $��]8���K�L\��Ki��q�d]t��q��Ki�L\���K��]8�$����w����پ�r��0���@:��fΌ�W��0郾\��eΌ�<:��&���}r����پw����x   x   �Im��!��/ُ� �����\�������!�/ُ��!���Im�_�P���3�#���u �(�׾�o���מ�᭍�>���vG��9���߭���מ��o��(�׾�u �!����3�e�P�x   x   �!��ߪ���؜��Ӥ�v���t����Ӥ��؜�ݪ���!���_j���K���-�������˾R��R����^���5���5���^��Y���R����˾�������-���K��_j�x   x   /ُ��؜�Y�lP������lP��W��؜�1ُ�b��� �a���A���#�PU��_�у��(����\�������v~������\��3���ك���_�LU���#���A� �a�f���x   x    ��Ӥ�lP��仱�滱�nP���Ӥ�!�È���;u��`T��X4�C��gw����ξ�����l������{��{�%����l��������ξlw��B���X4��`T��;u�È��x   x   ����v�������滱�����u��������m���!��g�c���B�=�#�R���߾빾-����A�z���r�=�z���-��#빾�߾T��:�#���B�]�c��!���m��x   x   \���t���lP��nP��u���\������䆿؉n��BN��.�������ž�$���-���z��wk��wk��z��-���$����ž�����.��BN�։n��䆿��x   x   �����Ӥ�W��Ӥ����������7t�XqU��6��6����� �о����`���u|���e�}e^���e�}u|��`�����)�о�����6���6�VqU�7t�!�����x   x   !𘿽؜��؜�!𘿺m���䆿7t�w�W��:������# پ����Q��0�~���a��S��S���a�2�~��Q�����  پ������:��W�7t��䆿�m��x   x   /ُ�ݪ��1ُ�È���!��؉n�XqU��:�����3�j�޾�ַ�����l���W_�MVK���D�KVK�W_�i��������ַ�i�޾�3�����:�YqU�׉n��!��ň��x   x   �!���!��b����;u�g�c��BN��6����3�kz��T������ȕ����]��UE�B,9�B,9��UE���]�ƕ�������T��fzྱ3����6��BN�b�c��;u�d���x   x   �Im��_j� �a��`T���B��.��6����j�޾�T���h���%���(]��{A�M1�}�+�M1��{A��(]��%���h���T��j�޾����6��.���B��`T� �a��_j�x   x   _�P���K���A��X4�=�#�������# پ�ַ������%��
�\���?�?/,���"���"�[/,���?��\��%�������ַ� پ������>�#��X4���A���K�g�P�x   x   ��3���-���#�C��R���� �о�������ȕ���(]���?���*����������*���?��(]�Ǖ���������,�о��P��>����#���-���3�6�x   x   #����PU�gw���߾��ž����Q��l�����]��{A�?/,�����������N/,�|A���]�m����Q�������ž�߾ow��MU���"���Q��Q�x   x   �u ����_⾥�ξ빾�$���`��0�~�W_��UE�M1���"������������"�`1��UE�W_�$�~��`���$��)빾��ξ�_⾎���u �H��d+�A��x   x   (�׾�˾у������-���-���u|���a�MVK�B,9�}�+���"�������"���+�<,9�OVK���a�yu|��-��-������Ӄ����˾)�׾I��<�E�F��x   x   �o��R��(����l�����z���e��S���D�B,9�M1�[/,���*�N/,�`1�<,9���D�ܨS���e��z� ���l��,���R���o��JR��+WľHƾ&WľGR��x   x   �מ�R����\�����A�z��wk�}e^��S�KVK��UE��{A���?���?�|A��UE�OVK�ܨS�oe^��wk�B�z�$����\��T����מ�aj��&����������&��jj��x   x   ᭍��^�������{���r��wk���e���a�W_���]��(]��\��(]���]�W_���a���e��wk�	�r��{������^��ޭ��(w��fJ�������WJ��1w��x   x   >����5���v~��{�=�z��z�}u|�2�~�i���ƕ���%���%��Ǖ��m���$�~�yu|��z�B�z��{��v~��5��:���X���j��.-��-!��.!��2-���j��W��x   x   vG���5������%������-���`���Q�����������h�����������Q���`���-�� ��$��������5��xG�����tG���������N:���������qG�����x   x   9����^���\���l��-���$���������ַ��T���T���ַ��������$��-���l���\���^��:������E1{��x�T[v�g�u�r�u�T[v��x�J1{����x   x   ߭��Y���3�������#빾��ž)�о  پi�޾fz�j�޾ پ,�о��ž)빾����,���T���ޭ��X��tG���x�^wr�oGo�@n�{Go�Uwr��x�mG��[��x   x   �מ�R��ك����ξ�߾�𾇊������3��3�����������߾��ξӃ��R���מ�(w���j������T[v�oGo��k���k�tGo�V[v� ����j��*w��x   x   �o����˾�_�lw��T�����6���������6���P��ow���_���˾�o��aj��fJ��.-�����g�u�@n���k��@n�j�u����0-��`J��hj��x   x   (�׾���LU�B��:�#��.���6��:��:��6��.�>�#�>��MU����)�׾JR��&���-!��N:��r�u�{Go�tGo�j�u�P:��.!���&��BR��x   x   �u �����#��X4���B��BN�VqU��W�YqU��BN���B��X4���#����u �I��+Wľ�������.!�����T[v�Uwr�V[v����.!���������-WľB��x   x   !����-���A��`T�]�c�։n�7t�7t�։n�b�c��`T���A���-�"��H��<�Hƾ�����2-�������x��x� ���0-�������CƾC�H��x   x   ��3���K� �a��;u��!���䆿!����䆿�!���;u� �a���K���3��Q�d+�E�&Wľ&��WJ���j��qG��J1{�mG���j��`J��&��-WľC�_+��Q�x   x   e�P��_j�f���È���m�������m��ň��d����_j�g�P�6��Q�A��F��GR��jj��1w��W��������[��*w��hj��BR��B��H���Q�6�x   x   �p�����M��R���$���$��R��K������p���!����d�`�A���!�N5���۾l���$�����8���9�������$��~l����۾P5���!�a�A��d��!��x   x   ���f\��2��`�ǿ�Eʿe�ǿ2��d\��������d���L\���8�f�������;�Ȭ������^����^�������Ȭ��;����l����8�L\�a������x   x   M��2��=Jʿ!�Ͽ"�Ͽ;Jʿ2��N����������;u��9O���+�����&�'���0���\���������\���0��'���&澬����+��9O��;u��������x   x   R��`�ǿ!�Ͽ�=ҿ!�Ͽa�ǿR���^������p��b�c�P>�������о옭��l���.��ـ���.���l��瘭��о�����P>�f�c��p������^��x   x   �$���Eʿ"�Ͽ!�Ͽ�Eʿ�$��M���cˠ�ԍ��~t��BN���*��x�����u��-����������������-���u�����~x���*��BN��~t�ԍ�bˠ�O���x   x   �$��e�ǿ;Jʿa�ǿ�$��g8���٤�D$��[B��u�Z��6�������Q�ƾ�$������2���v�2�������$��L�ƾ�������6�t�Z�`B��C$���٤�g8��x   x   R��2��2��R��M����٤�+����c��vb�R�>���r�;	Ҿ����s��J��m��m��I��s�����H	Ҿt���U�>�vb��c��,����٤�P���x   x   K��d\��N���^��cˠ�D$���c��%e�F`C��=#��3�{�ھ������� ��w"g�/�^��"g�� ��������t�ھ�3��=#�H`C�%e��c��@$��cˠ��^��x   x   �������������ԍ�[B��vb�F`C��%�*��fz��ַ�,��-����|b��RS��RS��|b����0���ַ�uz�1���%�B`C�	vb�_B��ԍ��������x   x   �p���������p���~t�u�Z�R�>��=#�*���m��T�������:����_���J��D���J���_��:�������T���m�*���=#�R�>�u�Z��~t��p��������x   x   �!��d����;u�b�c��BN��6����3�fz��T������ƕ����]��UE�B,9�B,9��UE���]�ȕ�������T��kzྫ3����6��BN�g�c��;u�b����!��x   x   ��d�L\��9O�P>���*����r�{�ھ�ַ�����ƕ���[]���B���2��t-���2���B��[]����������ַ���ھv������*�P>��9O�L\�w�d�Ccg�x   x   `�A���8���+����x����;	Ҿ���,���:����]���B�ߙ0���'��'�Ι0���B���]��:��=�����<	Ҿ���x������+���8�^�A�xF�xF�x   x   ��!�f�����������Q�ƾ������-�����_��UE���2���'�h�#��'��2��UE�q�_�)���������B�ƾ��⾃�����i��}�!��;'�/0)��;'�x   x   O5������&��о�u���$���s��� ���|b���J�B,9��t-��'��'� u-�8,9���J��|b�� ���s���$���u���о�&澍���U5���I.�N.���x   x   ��۾�;'��옭�-������J�w"g��RS��D�B,9���2�Ι0��2�8,9��D��RS�w"g�J�����-��ۘ��'��#�;��۾�c澞C�x�ﾪC��c�x   x   l���Ȭ��0���l�����2���m�/�^��RS���J��UE���B���B��UE���J��RS�7�^�(�m�9������l���0���Ȭ��l���O���ƾʾʾ�ƾ�O��x   x   �$�������\���.�������v��m��"g��|b���_���]��[]���]�q�_��|b�w"g�(�m��v������.���\�������$��Ơ���è�O��5��^���è�Ǡ��x   x   ����^�����ـ������2���I�� ������:��ȕ�������:��)���� ��J�9������׀������^�����詏�K钾{S����������zS��H钾婏�x   x   8��������.����������s�����0��������������=������s����������.������:���.郾�����f��� ��2:��� ���f������0郾x   x   9����^���\���l��-���$���������ַ��T���T���ַ��������$��-���l���\���^��:������E1{��x�T[v�g�u�r�u�T[v��x�J1{����x   x   ��������0��瘭��u��L�ƾH	Ҿt�ھuzྀm�kzྂ�ھ<	ҾB�ƾ�u��ۘ���0���������.郾E1{��q���k�!h�I�f�	!h���k� �q�P1{�/郾x   x   �$���Ȭ�'���о��⾚��t��3�1��*���3�v��������о'���Ȭ��$��詏������x���k��c�|�_�s�_��c���k��x�����⩏�x   x   ~l���;�&澈��~x�������=#��%��=#������x�����&�#�;�l��Ơ��K钾�f��T[v�!h�|�_�]�u�_�!h�W[v��f��K钾ʠ��x   x   ��۾�����������*��6�U�>�H`C�B`C�R�>��6���*�������������۾�O���è�{S��� ��g�u�I�f�s�_�u�_�G�f�o�u�� ��wS���è��O��x   x   P5�l����+�P>��BN�t�Z�vb�%e�	vb�u�Z��BN�P>���+�i��U5��c��ƾO������2:��r�u�	!h��c�!h�o�u�7:������b���ƾ�c�x   x   ��!���8��9O�f�c��~t�`B���c���c��_B���~t�g�c��9O���8�}�!����C�ʾ5������� ��T[v���k���k�W[v�� ������5��ʾ�C��x   x   a�A�L\��;u��p��ԍ�C$��,���@$��ԍ��p���;u�L\�^�A��;'�I.�x��ʾ^��zS���f���x� �q��x��f��wS��b��ʾ���J.��;'�x   x   �d�a���������bˠ��٤��٤�cˠ�������b���w�d�xF�/0)�N.��C��ƾ�è�H钾����J1{�P1{�����K钾�è��ƾ�C�J.�00)�xF�x   x   �!����������^��O���g8��P����^����������!��Ccg�xF��;'����c澈O��Ǡ��婏�0郾���/郾⩏�ʠ���O���c澔��;'�xF�=cg�x   x   ����xʿ,�׿Q�࿛{�O��-�׿�xʿ������/ُ�ju��L�%�'�J���ݾ(v���$��ݭ��Q���߭���$��'v����ݾJ� �'�ڍL�ou�2ُ����x   x   �xʿ��ڿ2}�����5}濑�ڿ�xʿi�������ň���Ki�ީ@�l��Bb��x�ξ�Ȭ�Y���_7��Z7��Y����Ȭ�v�ξHb��l���@��Ki�ƈ������k���x   x   ,�׿2}���l����6}�1�׿�Mſxׯ�����!��d�X� M1��N�Oy�'��.�����Q�����3���'��Ly��N��L1�`�X��!�����vׯ��Mſx   x   Q����l��m����N��>�Ͽga����ԍ�׉n���D�2��څ ��о������B㋾B㋾{�������оޅ �4����D�։n�ԍ���ea��@�Ͽx   x   �{������쿜{��$տ�¿nz���䖿_B��YqU��c.�������빾
����+��𷇾�+�����#빾��⾮���c.�YqU�^B���䖿nz���¿�$տx   x   O��5}�6}�N���$տ�3ſ>뱿���|���	vb��:��h������ž;���.A��������,A��<�����ž��� i��:�vb�}������=뱿�3ſ�$տx   x   -�׿��ڿ1�׿>�Ͽ�¿>뱿b������z�j�B`C����w�/�о%|��#��������,{�����$���|��)�оt����G`C�z�j����b���<뱿�¿@�Ͽx   x   �xʿ�xʿ�Mſga��nz��������O�m�`�G��%��3�( پ'K��BO���b���p��p��b��8O��+K��  پ�3��%�_�G�[�m�������nz��ba���Mſx   x   ���i���xׯ��󤿊䖿|���z�j�`�G���&�1��i�޾�������Ӏ�$�g�i�_�$�g�Ӏ��������i�޾1����&�`�G�z�j�|����䖿��xׯ�i���x   x   ����������ԍ�_B��	vb�B`C��%�1��uz��ַ�0������|b��RS��RS��|b�-���,���ַ�fz�*���%�F`C�vb�[B��ԍ�����������x   x   /ُ�ň���!��׉n�YqU��:�����3�i�޾�ַ�����i���W_�KVK���D�MVK�W_�l��������ַ�j�޾�3�����:�XqU�؉n��!��È��1ُ�ݪ��x   x   ju��Ki�d�X���D��c.��h�w�( پ���0��i���`Q^��eG��<��<��eG�qQ^�n���1����� پv� i��c.���D�^�X��Ki�pu�[7{�W7{�x   x   �L�ީ@� M1�2��������/�о'K���������W_��eG��'9�ym4��'9�
fG�W_�%������� K��,�о��󾶹�0���L1�ݩ@�ݍL�wT�)�V�lT�x   x   %�'�l���N�څ ������ž%|��BO��Ӏ��|b�KVK��<�ym4�fm4��<�MVK� }b�Ӏ�1O��!|����ž���ۅ ��N�i��'�'�0�/�:�3�;�3�0�/�x   x   J�Bb��Oy��о빾;���#����b��$�g��RS���D��<��'9��<���D��RS�+�g�c��"���/���)빾�оUy�Jb��J������$�����x   x   ��ݾx�ξ'������
���.A�������p�i�_��RS�MVK��eG�
fG�MVK��RS�{�_��p�����$A���������'��y�ξ��ݾ�<�Z�} ��l ��Z��<�x   x   (v���Ȭ�.������+������,{��p�$�g��|b�W_�qQ^�W_� }b�+�g��p��,{�����+�����,����Ȭ�$v��t���NjȾ
7;��ξ7;MjȾu���x   x   �$��Y�����B㋾𷇾��������b��Ӏ�-���l���n���%���Ӏ�c���������巇�P㋾��T����$��T��	,��V﫾MPN﫾	,��V��x   x   ݭ��_7��Q���B㋾�+��,A��$���8O������,������1������1O��"���$A���+��P㋾O���^7��ޭ��詏�Bϑ�V��������m������^���?ϑ�穏�x   x   Q���Z7����{�����<���|��*K������ַ��ַ���� K��!|��/�����������^7��K���X������9Ճ�����h��h������4Ճ�����\��x   x   ߭��Y���3�������#빾��ž)�о  پi�޾fz�j�޾ پ,�о��ž)빾����,���T���ޭ��X��tG���x�^wr�oGo�@n�{Go�Uwr��x�mG��[��x   x   �$���Ȭ�'���о��⾚��t��3�1��*���3�v��������о'���Ȭ��$��詏������x���k��c�|�_�s�_��c���k��x�����⩏�x   x   'v��v�ξLy�ޅ ���� i�����%���&��%���� i����ۅ �Uy�y�ξ$v��T��Bϑ�9Ճ�^wr��c�g�Z��X�|�Z�
�c�Pwr�5Ճ�Fϑ�Q��x   x   ��ݾHb���N�4���c.��:�G`C�^�G�`�G�F`C��:��c.�0���N�Jb����ݾt���	,��V�������oGo�|�_��X��X�x�_�oGo�����U���,��q���x   x   J�l���L1���D�YqU�vb�z�j�[�m�z�j�vb�XqU���D��L1�i��J��<�NjȾV﫾����h��@n�s�_�|�Z�x�_�u@n�h������T﫾LjȾ�<�x   x    �'��@�`�X�։n�^B��}���������|���[B��؉n�^�X�ݩ@�'�'���Z�
7;M�m��h��{Go��c�
�c�oGo�h���m��O
7;Z�
��x   x   ڍL��Ki��!��ԍ��䖿���b�������䖿ԍ��!���Ki�ݍL�0�/���} ����ξP��������Uwr���k�Pwr���������O��ξw ����3�/�x   x   ou�ƈ�������nz��=뱿<뱿nz���󤿫��È��pu�wT�:�3��$�l ��7;N﫾^���4Ճ��x��x�5Ճ�U���T﫾
7;w ���$�:�3�oT�x   x   2ُ�����vׯ�ea���¿�3ſ�¿ba��xׯ�����1ُ�[7{�)�V�;�3���Z�MjȾ	,��?ϑ�����mG������Fϑ�,��LjȾZ���:�3�0�V�\7{�x   x   ���k����Mſ@�Ͽ�$տ�$տ@�Ͽ�Mſi������ݪ��W7{�lT�0�/����<�u���V��穏�\��[��⩏�Q��q����<�
��3�/�oT�\7{�٪��x   x   r����' �	����( ���r�࿹xʿK��!𘿭q���jS�H++�h[	���ݾ|l���מ�O���J����מ�~l����ݾk[	�E++��jS��q�� �N���xʿx   x   ��z��j����k�x����~�ݿ�Mſ�^���m���q���D�n4�Vb��#�;R��f[�����e[��R���;Hb��v4���D��q��m���^���Mſ}�ݿx   x   ' �j�b�
�c�
�i�( ����6տba��cˠ��䆿�]�x!3��N��&�΃��[j��o���t���Vj��ك���&��N�x!3��]��䆿aˠ�ga���6տ��x   x   	�����c�
�������2��ۗ�v�ǿnz��@$��7t�y�F�4�������ξ-����V�����V��,�����ξ���4��z�F�7t�C$��oz��v�ǿ՗��2��x   x   ��k�i����u���濰�ϿN�������c���W��c.��x��߾$k�������x���x������'k���߾~x��c.�t�W��c�����M�����Ͽ���u��x   x   ( �x��( ��2�����bҿ�?��ˤ�����%e��:�������	þ%%���������%���	þ������:�%e����ˤ���?��cҿ���2��x   x   ������ۗ࿰�Ͽ�?��γ���s��[�m�H`C���~�����̾�M��k|���8���8��r|��N����̾������G`C�P�m��s��г���?����Ͽؗ���x   x   r��~�ݿ�6տv�ǿN���ˤ���s��afp�_�G��=#����%5Ծd߭��W��b���*$}�b����W��d߭�%5Ծ����=#�_�G�afp��s��ˤ��N���v�ǿ�6տ~�ݿx   x   �xʿ�Mſba��nz��������[�m�_�G��%��3�  پ+K��8O���b���p��p��b��BO��'K��( پ�3��%�`�G�O�m�������nz��ga���Mſ�xʿx   x   K���^��cˠ�@$���c��%e�H`C��=#��3�t�ھ������� ���"g�/�^�w"g�� ��������{�ھ�3��=#�F`C�%e��c��D$��cˠ��^��N��d\��x   x   !𘿹m���䆿7t��W��:������  پ����Q��2�~���a��S��S���a�0�~��Q�����# پ������:�w�W�7t��䆿�m��!𘿻؜��؜�x   x   �q���q��]�y�F��c.����~���%5Ծ+K�����2�~��*`��N��H�}N��*`��~����(K��%5Ծ��������c.�{�F��]��q��q���L�������L��x   x   �jS���D�x!3�4���x��𾔗̾d߭�8O��� ����a��N��CD��CD��N���a�� ��6O��d߭���̾��x�0��t!3���D��jS���]��:c��:c���]�x   x   H++�n4��N�����߾�	þ�M���W���b���"g��S��H��CD��H�ۨS�x"g��b���W��N���	þ�߾����N�u4�C++�h95�h�;��=�o�;�g95�x   x   h[	�Vb���&澪�ξ$k��%%��k|��b����p�/�^��S�}N��N�ۨS�6�^��p�\���v|��%%��)k����ξ�&�Jb��h[	�9�v��U��U��v��9�x   x   ��ݾ#�;΃��-����������8��*$}��p�w"g���a��*`���a�x"g��p�,$}�9�����������Ӄ��#�;��ݾ��љ��1���|	 �=���ԙ�����x   x   |l��R��[j���V���x������8��b����b��� ��0�~��~�� ���b��\���9������x���V��Jj��R���l��t����ɾ��ξ�Ҿ�Ҿ��ξ�ɾu���x   x   �מ�f[��o������x����r|���W��BO������Q�����6O���W��v|�����x����i���r[���מ�Ơ��	,��'�g��oD��g��'�
,��Ϡ��x   x   O������t����V������%��N��d߭�'K��������(K��d߭�N��%%�������V��i������O���(w��K钾V����s���ꔾ�ꔾ�s��U���I钾,w��x   x   J���e[��Vj��,���'k���	þ��̾%5Ծ( پ{�ھ# پ%5Ծ��̾�	þ)k�����Jj��r[��O���jΌ��j���f�������|��o+���|�������f���j��eΌ�x   x   �מ�R��ك����ξ�߾�𾇊������3��3�����������߾��ξӃ��R���מ�(w���j������T[v�oGo��k���k�tGo�V[v� ����j��*w��x   x   ~l���;�&澈��~x�������=#��%��=#������x�����&�#�;�l��Ơ��K钾�f��T[v�!h�|�_�]�u�_�!h�W[v��f��K钾ʠ��x   x   ��ݾHb���N�4���c.��:�G`C�^�G�`�G�F`C��:��c.�0���N�Jb����ݾt���	,��V�������oGo�|�_��X��X�x�_�oGo�����U���,��q���x   x   k[	�v4�x!3�z�F�t�W�%e�P�m�afp�O�m�%e�w�W�{�F�t!3�u4�h[	��뾠ɾ'��s���|���k�]��X�]�	�k��|���s��$��ɾ���x   x   E++���D��]�7t��c������s���s������c��7t��]���D�C++�9�љ����ξg���ꔾo+����k�u�_�x�_�	�k�m+���ꔾg����ξי��9�x   x   �jS��q��䆿C$�����ˤ��г��ˤ�����D$���䆿�q��jS�h95�v��1����ҾoD���ꔾ�|��tGo�!h�oGo��|���ꔾrD���Ҿ1���t��l95�x   x   �q���m��aˠ�oz��M����?���?��N���nz��cˠ��m���q����]�h�;�U��|	 ��Ҿg���s������V[v�W[v������s��g���Ҿ�	 �V��j�;���]�x   x    ��^��ga��v�ǿ��Ͽcҿ��Ͽv�ǿga���^��!��L���:c��=�U��=�����ξ'�U����f�� ����f��U���$���ξ1���V���=��:c��L��x   x   N���Mſ�6տ՗�����ؗ��6տ�MſN���؜������:c�o�;�v��ԙ���ɾ
,��I钾�j���j��K钾,���ɾי��t��j�;��:c������؜�x   x   �xʿ}�ݿ���2���u���2����~�ݿ�xʿd\���؜��L����]�g95�9����u���Ϡ��,w��eΌ�*w��ʠ��q������9�l95���]��L���؜�d\��x   x   �L�&��nb�g�pb�%���L���-�׿R������I���~�U�E++�J���۾�o���l��Rz���l���o����۾J�E++�{�U�H�������R��,�׿ ��x   x   &��&g�͈�͈�&g�'������@�ϿP�����d]t���D�l��������˾����T@��Z@��������˾����l����D�^]t���N���@�Ͽ����x   x   nb�͈���͈�ob�r�
�����ؗ��¿�٤�!����]��L1�����_�~��]����G��^���~���_⾬���L1��]�����٤��¿ח࿲���r�
�x   x   g�͈�͈�	g�Ȃ�ֈ���쿳�Ͽ<뱿,���7t���D���hw���s˾���������������s˾lw������D�7t�)���=뱿��Ͽ���׈�Ȃ�x   x   pb�&g�ob�Ȃ�<K����F�׿�?��b����c��VqU���*�Q��:�ھ�P���?���H���?���P��D�ھT����*�YqU��c��_����?��H�׿���;K�ǂ�x   x   %��'��r�
�ֈ����Y�ڿ���г�����vb���6������M���Ư��sp��wp��ǯ��W���������6�vb����ҳ�����O�ڿ���و�p�
�x   x   �L����������F�׿����ʦ��s��z�j�U�>��6�����SbƾF�����|ȍ���F���Sbƾ�����6�U�>�z�j��s���ʦ����F�׿��쿯�����x   x   ����ؗ࿳�Ͽ�?��г���s��P�m�G`C���������̾N��r|���8���8��k|���M����̾~�����H`C�[�m��s��γ���?����Ͽۗ�����x   x   -�׿@�Ͽ�¿<뱿b������z�j�G`C����t�)�о|��$��������,{�����#���%|��/�оw����B`C�z�j����b���>뱿�¿>�Ͽ1�׿��ڿx   x   R��P����٤�,����c��vb�U�>���t�H	Ҿ����s���I��m��m�J��s�����;	Ҿr���R�>�vb��c��+����٤�M���R��2��2��x   x   ������!���7t�VqU���6��6�����)�о����`��}u|���e�}e^���e��u|��`����� �о�����6��6�XqU�7t������ ����Ӥ�W��Ӥ�x   x   I���d]t��]���D���*���������̾|���s��}u|�N@c�7�V�L�V�=@c��u|��s��|����̾��������*���D��]�c]t�F���'-����������'-��x   x   ~�U���D��L1���Q�����SbƾN��$����I���e�7�V���Q�>�V���e�J�(���N��Rbƾx��P������L1���D�x�U���b�P3k�on�B3k���b�x   x   E++�l�����hw��:�ھM���F���r|�������m�}e^�L�V�>�V�ve^��m�����q|��@���J���D�ھow�����i��C++�L7�O�?�*D�(D�M�?�M7�x   x   J������_⾐s˾�P��Ư�����8���,{��m���e�=@c���e��m��,{��8���𓾹����P���s˾�_⾍���J�9�Y������� ����Z��9�x   x   ��۾��˾~������?��sp��|ȍ��8������J��u|��u|�J������8��vȍ�np���?�����~����˾��۾�<�љ������"��"����ݙ���<�x   x   �o������]��������H��wp����k|��#����s���`���s��(���q|����np���H������i��������o���O��NjȾ��ξ?.Ӿ��Ծ;.Ӿ��ξQjȾ�O��x   x   �l��T@���G�������?��ǯ��F����M��%|��������|��N��@��������?�������G��^@���l��aj���è�V﫾g��d���g��� g��N﫾�è�lj��x   x   Rz��Z@��^�������P��W���Sbƾ��̾.�о;	Ҿ �о��̾RbƾJ����P�����i���^@��Lz��;:��fJ��{S�������ꔾ픾�ꔾ����yS��[J��=:��x   x   �l������~���s˾D�ھ�������~���w�r���������x��D�ھ�s˾~�������l��;:��n-��.-��� ��h��o+��r+��h��� ��2-��q-��<:��x   x   �o����˾�_�lw��T�����6���������6���P��ow���_���˾�o��aj��fJ��.-�����g�u�@n���k��@n�j�u����0-��`J��hj��x   x   ��۾�����������*��6�U�>�H`C�B`C�R�>��6���*�������������۾�O���è�{S��� ��g�u�I�f�s�_�u�_�G�f�o�u�� ��wS���è��O��x   x   J�l���L1���D�YqU�vb�z�j�[�m�z�j�vb�XqU���D��L1�i��J��<�NjȾV﫾����h��@n�s�_�|�Z�x�_�u@n�h������T﫾LjȾ�<�x   x   E++���D��]�7t��c������s���s������c��7t��]���D�C++�9�љ����ξg���ꔾo+����k�u�_�x�_�	�k�m+���ꔾg����ξי��9�x   x   {�U�^]t����)���_���ҳ���ʦ�γ��b���+������b]t�x�U�K7�Y�����?.Ӿd���픾r+���@n�G�f�u@n�m+��픾_���7.Ӿ���_��N7�x   x   H������٤�=뱿�?���������?��>뱿�٤���F�����b�O�?�����"���Ծg����ꔾh��j�u�o�u�h���ꔾ_�����Ծ�"����L�?���b�x   x   ����N����¿��ϿH�׿O�ڿF�׿��Ͽ�¿M�������'-��P3k�*D��� ��"�;.Ӿ g������� ������ ������g��7.Ӿ�"��� �+D�L3k�(-��x   x   R��@�Ͽח࿍�쿫���򿏫�ۗ�>�ϿR���Ӥ�����on�(D���������ξN﫾yS��2-��0-��wS��T﫾��ξ������+D�gn������Ӥ�x   x   ,�׿�쿲���׈�;K�و�������1�׿2��W�����B3k�M�?�Z��ݙ��QjȾ�è�[J��q-��`J���è�LjȾי��_��L�?�L3k�����Y�2��x   x    ����r�
�Ȃ�ǂ�p�
������ڿ2���Ӥ�'-����b�M7�9��<꾃O��lj��=:��<:��hj���O���<�9�N7���b�(-���Ӥ�2����ڿx   x   ����:#���'���'��:#����%��( �O�࿨$��\���F����jS�%�'�R5�2�׾@ط�f5��`5��Bط�(�׾P5� �'��jS�H���\����$��L��' �&��x   x   �:#�*�},� *��:#�uw�p�
��2���$տg8�����q�ک@�d������`ɾ���f
������`ɾ���l���@��q���e8���$տ�2��s�
�sw�x   x   ��'�},�},���'�n�� h�و��濂3ſ�٤��䆿b�X���+�OU��ܾڌ��t��t��،��دܾLU���+�`�X��䆿�٤��3ſ��ֈ�h�o��x   x   ��'� *���'�!�aj�������cҿ=뱿C$��։n�P>�>��&���@Ǿa@���\��`@���@Ǿ1��B��P>�։n�C$��=뱿cҿ�����`j�!�x   x   �:#��:#�n��aj�I�
�!w��O�ڿ�?�����`B���BN�=�#�(��\Ӿ����社	褾����\Ӿ(�:�#��BN�^B������?��R�ڿ!w��H�
�bj�o��x   x   ���uw� h����!w��D�ݿ���ˤ��}���t�Z��.���
���޾����̣������̣������޾��
��.�t�Z�}���ˤ�����D�ݿ!w����� h�uw�x   x   %��p�
�و����O�ڿ���ҳ�����vb��6������W���ǯ��wp��sp��Ư��M����������6�vb����г�����Y�ڿ���ֈ�r�
�'��x   x   ( ��2����cҿ�?��ˤ�����%e��:�������	þ%���������%%���	þ������:�%e����ˤ���?���bҿ���2��( �x��x   x   O���$տ�3ſ=뱿���}���vb��:� i������ž<���,A��������.A��;�����ž����h��:�	vb�|������>뱿�3ſ�$տN��6}�5}�x   x   �$��g8���٤�C$��`B��t�Z��6�������L�ƾ�$������2���v�2�������$��Q�ƾ�������6�u�Z�[B��D$���٤�g8���$��a�ǿ;Jʿe�ǿx   x   \������䆿։n��BN��.�������ž�$���-���z��wk��wk��z��-���$����ž�����.��BN�؉n��䆿��\���u���nP��lP��t���x   x   F����q�b�X�P>�=�#���
�����	þ<��������z���g��a���g�#�z�����5����	þ~�边�
�>�#�P>�^�X��q�F����؋���쒿���؋�x   x   �jS�ک@���+�>��(���޾W���%��,A��2���wk��a���a��wk�(��$A��%��R�����޾(�>����+�ݩ@��jS���b���m���s�ʭs���m���b�x   x   %�'�d��OU�&���\Ӿ���ǯ��������v��wk���g��wk���v������ɯ������\Ӿ!��MU�i��'�'�h95�O�?��2F��tH��2F�S�?�h95�x   x   R5�����ܾ�@Ǿ����̣�wp��������2���z�#�z�(��������rp���̣�����@Ǿ�ܾ���U5���v�����z6"�w6"����z����x   x   2�׾�`ɾڌ��a@���社����sp����.A�������-������$A����rp������褾[@��挻��`ɾ)�׾�c�Z�1����"��F��"�,���&Z��c�x   x   @ط����t���\��	褾�̣�Ư��%%��;����$���$��5���%��ɯ���̣�褾�\��)t�����:ط�JR���ƾ
7;�Ҿ��Ծ��Ծ�Ҿ7;�ƾ?R��x   x   f5��f
��t��`@��������M����	þ��žQ�ƾ��ž�	þR���������[@��)t��`
��\5��*���&��O��MoD��g���cD��SZ��&��$���x   x   `5�����،���@Ǿ�\Ӿ��޾��辟������~����޾�\Ӿ�@Ǿ挻����\5���<��,��������m���ꔾ�ꔾ�m�������,���<��x   x   Bط��`ɾدܾ1��(���
�������h��������
�(�!���ܾ�`ɾ:ط�*���,���[��-!��2:��h���|��h��0:��/!���[��,��&���x   x   (�׾���LU�B��:�#��.���6��:��:��6��.�>�#�>��MU����)�׾JR��&���-!��N:��r�u�{Go�tGo�j�u�P:��.!���&��BR��x   x   P5�l����+�P>��BN�t�Z�vb�%e�	vb�u�Z��BN�P>���+�i��U5��c��ƾO������2:��r�u�	!h��c�!h�o�u�7:������b���ƾ�c�x   x    �'��@�`�X�։n�^B��}���������|���[B��؉n�^�X�ݩ@�'�'���Z�
7;M�m��h��{Go��c�
�c�oGo�h���m��O
7;Z�
��x   x   �jS��q��䆿C$�����ˤ��г��ˤ�����D$���䆿�q��jS�h95�v��1����ҾoD���ꔾ�|��tGo�!h�oGo��|���ꔾrD���Ҿ1���t��l95�x   x   H������٤�=뱿�?���������?��>뱿�٤���F�����b�O�?�����"���Ծg����ꔾh��j�u�o�u�h���ꔾ_�����Ծ�"����L�?���b�x   x   \���e8���3ſcҿR�ڿD�ݿY�ڿ�bҿ�3ſg8��\����؋���m��2F�z6"��F���ԾcD���m��0:��P:��7:���m��rD����Ծ�F�x6"��2F���m��؋�x   x   �$���$տ�濪��!w��!w��������$տ�$��u�������s��tH�w6"��"��ҾS����/!��.!������O�Ҿ�"�x6"��tH�ɭs���t���x   x   L���2��ֈ����H�
����ֈ��2��N��a�ǿnP��쒿ʭs��2F����,���7;Z����[���b��
7;1�������2F�ɭs�쒿nP��`�ǿx   x   ' �s�
�h�`j�bj� h�r�
�( �6}�;JʿlP������m�S�?�z��&Z��ƾ&��,��,��&���ƾZ�t��L�?���m���nP��;Jʿ6}�x   x   &��sw�o��!�o��uw�'��x��5}�e�ǿt����؋���b�h95����c�?R��$����<��&���BR���c�
��l95���b��؋�t���`�ǿ6}�|��x   x   -�.�~k6��9�k6�-�.��:#�pb����{㿪$�������q���L���!��u �@`Ӿ�&��R����&��F`Ӿ�u ���!�ڍL��q�������$���{���mb��:#�x   x   ~k6�m�;�n�;�k6��,�o��ǂ��u���$տO����m���Ki���8������$�ƾ,��5��%�ƾ�������8��Ki��m��N����$տ�u��Ȃ�n���,�x   x   �9�n�;��9��_1��~%�bj�;K����¿cˠ��!���9O���#�u�B�վ�D�������D��B�վw���#��9O��!��aˠ��¿��;K�`j��~%��_1�x   x   k6�k6��_1���'�Ս�H�
���򿶯Ͽnz��ԍ�]�c��X4� ��澓�¾ñ��±���¾� ���X4�f�c�ԍ�oz����Ͽ���J�
�Ս���'��_1�x   x   -�.��,��~%�Ս�A��!w��H�׿M����䖿�~t���B��5�=���%˾�j���M���j��%˾=����5���B��~t��䖿M���H�׿!w��A��Ս��~%��,�x   x   �:#�o��bj�H�
�!w��R�ڿ�?�����^B���BN�:�#�(��\Ӿ���	褾�社����\Ӿ(�=�#��BN�`B������?��O�ڿ!w��I�
�aj�n���:#�x   x   pb�ǂ�;K����H�׿�?��_����c��YqU���*�T��D�ھ�P���?���H���?���P��:�ھQ����*�VqU��c��b����?��F�׿���<K�Ȃ�ob�&g�x   x   ���u���濶�ϿM�������c��t�W��c.�~x��߾'k�������x���x������$k���߾�x��c.��W��c�����N�����Ͽ���u����i�k�x   x   �{��$տ�¿nz���䖿^B��YqU��c.�������#빾����+��𷇾�+��
���빾��⾰���c.�YqU�_B���䖿nz���¿�$տ�{�������x   x   �$��O���cˠ�ԍ��~t��BN���*�~x�����u��-����������������-���u����⾀x���*��BN��~t�ԍ�cˠ�M����$���Eʿ!�Ͽ"�Ͽ�Eʿx   x   �����m���!��]�c���B�:�#�T���߾#빾-����=�z���r�A�z���-��빾�߾R��=�#���B�g�c��!���m�� ���u�������滱�����v���x   x   �q���Ki��9O��X4��5�(�D�ھ'k��������=�z���m���m�E�z�������2k��A�ھ(��5��X4��9O��Ki��q��'-����1���6�����$-��x   x   �L���8���#� ��=����\Ӿ�P�������+��������r���m���r������+�������P���\Ӿ0���!����#���8�ݍL���]�P3k���s�F�v���s�H3k���]�x   x   ��!���u��%˾����?���x��𷇾����A�z�E�z�������x���?�����%˾��x���}�!�0�/�h�;�*D��tH��tH�(D�h�;�1�/�x   x   �u ����B�վ��¾�j��	褾�H���x���+�����������+���x���H��	褾�j����¾A�վ����u �����U���� �w6"��� �Q������x   x   @`Ӿ$�ƾ�D��ñ��M���社�?������
���-��-����������?��	褾�M���±��D���ƾQ`ӾI�ྞC�} ��|	 ��"��"��	 �r ���C�H��x   x   �&��,�������±��j������P��$k��빾�u��빾2k���P������j���±�����'���&���r��+Wľʾ��ξ�Ҿ;.Ӿ�Ҿ��ξʾ3Wľyr��x   x   R���5���D����¾%˾�\Ӿ:�ھ�߾�������߾A�ھ�\Ӿ%˾��¾�D��'��`���qޭ�®������5��Pg�� g��S5������̮��iޭ�x   x   �&��%�ƾB�վ�=���(�Q���x�����x�R��(�0�����A�վ�ƾ�&��qޭ��椾�=��������������s��������������=���椾gޭ�x   x   F`Ӿ���w� ���5�=�#���*��c.��c.���*�=�#��5�!��x����Q`Ӿ�r��®���=����.!��� ����������� ��/!�����=��̮��}r��x   x   �u �����#��X4���B��BN�VqU��W�YqU��BN���B��X4���#����u �I��+Wľ�������.!�����T[v�Uwr�V[v����.!���������-WľB��x   x   ��!���8��9O�f�c��~t�`B���c���c��_B���~t�g�c��9O���8�}�!����C�ʾ5������� ��T[v���k���k�W[v�� ������5��ʾ�C��x   x   ڍL��Ki��!��ԍ��䖿���b�������䖿ԍ��!���Ki�ݍL�0�/���} ����ξP��������Uwr���k�Pwr���������O��ξw ����3�/�x   x   �q���m��aˠ�oz��M����?���?��N���nz��cˠ��m���q����]�h�;�U��|	 ��Ҿg���s������V[v�W[v������s��g���Ҿ�	 �V��j�;���]�x   x   ����N����¿��ϿH�׿O�ڿF�׿��Ͽ�¿M�������'-��P3k�*D��� ��"�;.Ӿ g������� ������ ������g��7.Ӿ�"��� �+D�L3k�(-��x   x   �$���$տ�濪��!w��!w��������$տ�$��u�������s��tH�w6"��"��ҾS����/!��.!������O�Ҿ�"�x6"��tH�ɭs���t���x   x   �{��u��;K�J�
�A��I�
�<K��u���{��Eʿ����1���F�v��tH��� ��	 ���ξ5����������5����ξ�	 ��� ��tH�7�v�3��������Eʿx   x   ��Ȃ�`j�Ս�Ս�aj�Ȃ�����!�Ͽ滱�6�����s�(D�Q��r ��ʾ�����=���=������ʾw ��V��+D�ɭs�3���仱� �Ͽ��x   x   mb�n���~%���'��~%�n��ob�i���"�Ͽ������H3k�h�;����C�3Wľ̮���椾̮��-Wľ�C���j�;�L3k������� �Ͽ��j�x   x   �:#��,��_1��_1��,��:#�&g�k����Eʿv���$-����]�1�/���H��yr��iޭ�gޭ�}r��B�ྔ�3�/���]�(-��t����Eʿ��j�&g�x   x   A�V�F�W�F�A�k6���'�g�	��Q��R�� �nu�\�A�#���$��f�ξ�绾�绾`�ξ�$��!��a�A�ou� �R��L����	g���'�k6�x   x   V�F��I�U�F�ZX>��_1�!�Ȃ��2��@�Ͽ�^��È��L\���-���	�<5�3�ľN4��4�ľ35���	���-�L\�ƈ���^��@�Ͽ�2��Ȃ�!��_1�[X>�x   x   W�F�U�F�aA�rl6���'�`j�׈�՗�ea������;u���A����y����ξ=��=����ξ�x�������A��;u����ga��ח�ֈ�`j���'�pl6�aA�x   x   A�ZX>�rl6�� *�Ս�������v�ǿ�󤿍p���`T���'�2�}^ھ�ﾾ�����ﾾ}^ھ2���'��`T��p����v�ǿ��쿪��Ս�� *�rl6�ZX>�x   x   k6��_1���'�Ս�J�
���򿯯Ͽoz��ԍ�f�c��X4� ��澖�¾�±�ñ���¾� ���X4�]�c�ԍ�nz����Ͽ���H�
�Ս���'��_1�k6�x   x   ��'�!�`j�������cҿ=뱿C$��։n�P>�B��1���@Ǿ`@���\��a@���@Ǿ&��>��P>�։n�C$��=뱿cҿ�����aj�!���'� *�x   x   g�Ȃ�׈���쿯�Ͽ=뱿)���7t���D���lw���s˾���������������s˾hw������D�7t�,���<뱿��Ͽ���ֈ�Ȃ�	g�͈�͈�x   x   	���2��՗�v�ǿoz��C$��7t�z�F�4�������ξ,����V�����V��-�����ξ���4��y�F�7t�@$��nz��v�ǿۗ��2�������c�
����x   x   Q��@�Ͽea����ԍ�։n���D�4��ޅ ��о����{��B㋾B㋾�������оڅ �2����D�׉n�ԍ���ga��>�ϿN����m��l����x   x   R���^������p��f�c�P>�������о瘭��l���.��ـ���.���l��옭��о�����P>�b�c��p������^��R��a�ǿ!�Ͽ�=ҿ!�Ͽ`�ǿx   x    �È���;u��`T��X4�B��lw����ξ�����l��%����{��{�����l��������ξgw��C���X4��`T��;u�È��!��Ӥ�nP��滱�仱�lP���Ӥ�x   x   nu�L\���A���'� ��1��s˾,���{���.���{���u�!�{��.�����'����s˾+������'���A�L\�pu��L������쒿6���쒿�����L��x   x   \�A���-����2���@Ǿ����V��B㋾ـ���{�!�{�΀��G㋾�V������@Ǿ��7������-�^�A�wT��:c�on�ʭs���s�rn��:c�tT�x   x   #����	�y��}^ھ��¾`@��������B㋾�.������.��G㋾�򓾯���`@����¾�^ھ�x����	�"���;'�:�3��=�(D��2F�(D�#�=�9�3��;'�x   x   �$��<5ᾈ�ξ�ﾾ�±��\�������V�����l���l������V�������\���±��ﾾ��ξ@5ᾣ$��H��I.��$�U��������Q���$�L.�F��x   x   f�ξ3�ľ=������ñ�a@�����-�������옭�����'������`@���±�����	=��8�ľk�ξ��پ<�x��l ��=������,���r ��{��?循�پx   x   �绾N4��=���ﾾ��¾�@Ǿ�s˾��ξ�о�о��ξ�s˾�@Ǿ��¾�ﾾ	=��T4���绾I��C���Hƾʾ7;��ξ��ξ7;ʾ>ƾI���1I��x   x   �绾4�ľ��ξ}^ھ�&��hw�����څ ����gw��+���澆^ھ��ξ8�ľ�绾hX���а��������^��N﫾'�N﫾Z����������а�uX��x   x   `�ξ35��x��2� ��>����4��2����C����7��x��@5�k�ξI���а��(���=���zS��^���U���yS����=���(���а�3I��x   x   �$����	������'��X4�P>���D�y�F���D�P>��X4���'������	��$����پC�������=���[��2-���f��4Ճ��f��2-���[���=�����H�����پx   x   !����-���A��`T�]�c�։n�7t�7t�׉n�b�c��`T���A���-�"��H��<�Hƾ�����2-�������x��x� ���0-�������CƾC�H��x   x   a�A�L\��;u��p��ԍ�C$��,���@$��ԍ��p���;u�L\�^�A��;'�I.�x��ʾ^��zS���f���x� �q��x��f��wS��b��ʾ���J.��;'�x   x   ou�ƈ�������nz��=뱿<뱿nz���󤿫��È��pu�wT�:�3��$�l ��7;N﫾^���4Ճ��x��x�5Ճ�U���T﫾
7;w ���$�:�3�oT�x   x    ��^��ga��v�ǿ��Ͽcҿ��Ͽv�ǿga���^��!��L���:c��=�U��=�����ξ'�U����f�� ����f��U���$���ξ1���V���=��:c��L��x   x   R��@�Ͽח࿍�쿫���򿏫�ۗ�>�ϿR���Ӥ�����on�(D���������ξN﫾yS��2-��0-��wS��T﫾��ξ������+D�gn������Ӥ�x   x   L���2��ֈ����H�
����ֈ��2��N��a�ǿnP��쒿ʭs��2F����,���7;Z����[���b��
7;1�������2F�ɭs�쒿nP��`�ǿx   x   ��Ȃ�`j�Ս�Ս�aj�Ȃ�����!�Ͽ滱�6�����s�(D�Q��r ��ʾ�����=���=������ʾw ��V��+D�ɭs�3���仱� �Ͽ��x   x   	g�!���'�� *���'�!�	g����m���=ҿ仱�쒿rn�#�=��$�{��>ƾ����(�����Cƾ����$��=�gn�쒿仱��=ҿm�����x   x   ��'��_1�pl6�rl6��_1���'�͈�c�
�l��!�ϿlP�������:c�9�3�L.�?�I����а��а�H���C�J.�:�3��:c�����nP�� �Ͽm��c�
�̈�x   x   k6�[X>�aA�ZX>�k6� *�͈������`�ǿ�Ӥ��L��tT��;'�F����پ1I��uX��3I����پH���;'�oT��L���Ӥ�`�ǿ�����̈� *�x   x   p�O�h�R�r�O�W�F��9���'�nb�' �,�׿M��/ُ�y�d���3��R�q`��Wʾ�����Wʾm`辀R���3��d�2ُ�N��,�׿' �mb���'��9�W�F�x   x   h�R�h�R���L�aA��_1�o��r�
��쿟Mſ����f�����K��> �V? �q׾��þ��þq׾Z? ��> ���K�a��������Mſ��s�
�n���_1�`A���L�x   x   r�O���L�_�C�pl6��~%�h������6տvׯ���� �a���1�����#�ɏȾA���ɏȾ�#������1� �a����vׯ��6տ����h��~%�pl6�_�C���L�x   x   W�F�aA�pl6���'�`j�ֈ�ח�ga������;u���A�����x����ξ=��=����ξy�������A��;u����ea��՗�׈�`j���'�rl6�aA�U�F�x   x   �9��_1��~%�`j�;K����¿aˠ��!���9O���#�w�B�վ�D�������D��B�վu���#��9O��!��cˠ��¿��;K�bj��~%��_1��9�n�;�x   x   ��'�o��h�ֈ��濇3ſ�٤��䆿`�X���+�LU�دܾ،��t��t��ڌ���ܾOU���+�b�X��䆿�٤��3ſ��و� h�n����'�},�},�x   x   nb�r�
�����ח��¿�٤�����]��L1�����_�~��^����G��]���~���_⾬���L1��]�!����٤��¿ؗ࿯���r�
�ob�͈���͈�x   x   ' ����6տga��aˠ��䆿�]�x!3��N��&�ك��Vj��t���o���[j��΃���&��N�x!3��]��䆿cˠ�ba���6տ��( �i�c�
�b�
�j�x   x   ,�׿�Mſvׯ�����!��`�X��L1��N�Ly�'��3�����Q�����.���'��Oy��N� M1�d�X��!�����xׯ��Mſ1�׿6}���l����2}�x   x   M����������;u��9O���+�����&�'���0���\���������\���0��'���&澫����+��9O��;u��������N��2��;Jʿ"�Ͽ!�Ͽ=Jʿ2��x   x   /ُ�f��� �a���A���#�LU��_�ك��3����\�������v~������\��(���у���_�PU���#���A� �a�b���1ُ��؜�W�lP������lP��Y��؜�x   x   y�d���K���1����w�دܾ~��Vj��������v~��v~������Hj��~��ܾ߯v������1���K�w�d�[7{���������������������\7{�x   x   ��3��> �����x��B�վ،��^���t���Q�������������N���h���e���茻�F�վy������> ���3�xF�)�V��:c�B3k���m�H3k��:c�!�V�xF�x   x   �R�V? ��#澇�ξ�D��t���G��o������\���\����h����G��&t���D����ξ�#�U? ��R��Q�/0)�;�3�o�;�M�?�S�?�h�;�9�3�10)��Q�x   x   q`�q׾ɏȾ=������t��]���[j��.����0��(���Hj��e���&t������=��Ⱦ	q׾f`�w��d+�N.���v��Z��z����L.�b+�w��x   x   �Wʾ��þA���=���D��ڌ��~��΃��'��'��у��~��茻��D��=��=�����þ�Wʾ�ҾJ�۾E循C�Z�ԙ��ݙ��&Z�C�?�;�۾�Ҿx   x   ������þɏȾ��ξB�վ�ܾ�_⾝&�Oy群&澐_�ܾ߯F�վ��ξȾ��þ����s���
��J���&Wľ�ƾMjȾ�ɾQjȾ�ƾ3WľI����
��s��x   x   �Wʾq׾�#�y��u�OU�����N��N����PU�v�y���#�	q׾�Wʾs�������а�Ǯ��&���è�	,��
,���è�&��̮���а�����s��x   x   m`�Z? ���������#���+��L1�x!3� M1���+���#�������U? �f`��Ҿ�
���а��椾,��WJ��H钾?ϑ�I钾[J��,���椾�а��
���Ҿx   x   �R��> ���1���A��9O�b�X��]��]�d�X��9O���A���1��> ��R�w��J�۾J���Ǯ��,��j-���j�����������j��q-��,��̮��H���2�۾w��x   x   ��3���K� �a��;u��!���䆿!����䆿�!���;u� �a���K���3��Q�d+�E�&Wľ&��WJ���j��qG��J1{�mG���j��`J��&��-WľC�_+��Q�x   x   �d�a���������bˠ��٤��٤�cˠ�������b���w�d�xF�/0)�N.��C��ƾ�è�H钾����J1{�P1{�����K钾�è��ƾ�C�J.�00)�xF�x   x   2ُ�����vׯ�ea���¿�3ſ�¿ba��xׯ�����1ُ�[7{�)�V�;�3���Z�MjȾ	,��?ϑ�����mG������Fϑ�,��LjȾZ���:�3�0�V�\7{�x   x   N���Mſ�6տ՗�����ؗ��6տ�MſN���؜������:c�o�;�v��ԙ���ɾ
,��I钾�j���j��K钾,���ɾי��t��j�;��:c������؜�x   x   ,�׿�쿲���׈�;K�و�������1�׿2��W�����B3k�M�?�Z��ݙ��QjȾ�è�[J��q-��`J���è�LjȾי��_��L�?�L3k�����Y�2��x   x   ' �s�
�h�`j�bj� h�r�
�( �6}�;JʿlP������m�S�?�z��&Z��ƾ&��,��,��&���ƾZ�t��L�?���m���nP��;Jʿ6}�x   x   mb�n���~%���'��~%�n��ob�i���"�Ͽ������H3k�h�;����C�3Wľ̮���椾̮��-Wľ�C���j�;�L3k������� �Ͽ��j�x   x   ��'��_1�pl6�rl6��_1���'�͈�c�
�l��!�ϿlP�������:c�9�3�L.�?�I����а��а�H���C�J.�:�3��:c�����nP�� �Ͽm��c�
�̈�x   x   �9�`A�_�C�aA��9�},���b�
���=JʿY�����!�V�10)�b+�;�۾�
�������
��2�۾_+�00)�0�V�����Y�;Jʿ��c�
���},�x   x   W�F���L���L�U�F�n�;�},�͈�j�2}�2���؜�\7{�xF��Q�w���Ҿs��s���Ҿw���Q�xF�\7{��؜�2��6}�j�̈�},�m�;�x   x   qMY�pMY�h�R�V�F�~k6��:#�&����xʿ����!��^�P�$�r�&�۾�Ǿ�Ǿ#�۾q�$�e�P��!������xʿ ��&���:#�k6�W�F�g�R�x   x   pMY���U���L�[X>��,�sw���}�ݿk�������_j��]8������Y�ξ��ľY�ξ������]8��_j����k���}�ݿ��sw��,�[X>���L���U�x   x   h�R���L�`A��_1�n��s�
��쿜Mſ����a�����K��> �Z? �q׾��þ��þq׾V? ��> ���K�f��������Mſ��r�
�o���_1�aA���L�h�R�x   x   V�F�[X>��_1�!�Ȃ��2��@�Ͽ�^��ƈ��L\���-���	�35�4�ľN4��3�ľ<5���	���-�L\�È���^��@�Ͽ�2��Ȃ�!��_1�ZX>�U�F��I�x   x   ~k6��,�n��Ȃ��u���$տN����m���Ki���8������%�ƾ5��,��$�ƾ�������8��Ki��m��O����$տ�u��ǂ�o���,�k6�n�;�m�;�x   x   �:#�sw�s�
��2���$տe8�����q��@�l������`ɾ���f
������`ɾ���d��ک@��q���g8���$տ�2��p�
�uw��:#� *�},�*�x   x   &������@�ϿN�����^]t���D�l��������˾����Z@��T@��������˾����l����D�d]t���P���@�Ͽ����'��&g�͈�͈�&g�x   x   ��}�ݿ�Mſ�^���m���q���D�v4�Hb���;R��e[�����f[��R��#�;Vb��n4���D��q��m���^���Mſ~�ݿ��x��k����j�z��x   x   �xʿk�������ƈ���Ki��@�l��Hb��v�ξ�Ȭ�Y���Z7��_7��Y����Ȭ�x�ξBb��l��ީ@��Ki�ň������i����xʿ��ڿ5}�����2}濐�ڿx   x   ������a���L\���8�l�������;�Ȭ������^����^�������Ȭ��;����f����8�L\�d���������d\��2��e�ǿ�Eʿ`�ǿ2��f\��x   x   �!���_j���K���-��������˾R��Y����^���5���5���^��R���R���˾�������-���K��_j��!��ݪ���؜��Ӥ�t���v����Ӥ��؜�ߪ��x   x   ^�P��]8��> ���	�����`ɾ����e[��Z7����5���[7��p[�������`ɾ����	��> ��]8�g�P�Ccg�W7{��L��'-���؋�$-���L��\7{�Hcg�x   x   $���Z? �35�%�ƾ���Z@�����_7���^���^��[7�����e@������ƾ;5�W? �!��$�6�xF�lT���]���b���b���]�tT�xF�6�x   x   r����q׾4�ľ5��f
��T@��f[��Y�������R���p[��e@��b
��"��2�ľq׾���u�����Q��;'�0�/�g95�M7�h95�1�/��;'��Q����x   x   &�۾Y�ξ��þN4��,���������R���Ȭ��Ȭ�R���������"��U4����þ`�ξ%�۾���w��A������9�9�����F��w�����x   x   �Ǿ��ľ��þ3�ľ$�ƾ�`ɾ��˾#�;x�ξ�;�˾�`ɾ�ƾ2�ľ��þȠľ�Ǿ3V̾�Ҿ��پF���c��<�����<��c�H�ྪ�پ�Ҿ(V̾x   x   �ǾY�ξq׾<5���꾑�����Vb��Bb������������;5�q׾`�ξ�ǾC{¾s��I���r��GR���O��u���u����O��?R��yr��1I��s��={¾x   x   #�۾���V? ���	���d��l��n4�l��f�����	�W? ����%�۾3V̾s��fX��jޭ�0���jj��Ǡ��V��Ϡ��lj��$���iޭ�uX��s��-V̾x   x   q����> ���-���8�ک@���D���D�ީ@���8���-��> �!��u�����ҾI��jޭ��<��@:��1w��婏�穏�,w��=:���<��gޭ�3I���Ҿ���x   x   $��]8���K�L\��Ki��q�d]t��q��Ki�L\���K��]8�$����w����پ�r��0���@:��fΌ�W��0郾\��eΌ�<:��&���}r����پw����x   x   e�P��_j�f���È���m�������m��ň��d����_j�g�P�6��Q�A��F��GR��jj��1w��W��������[��*w��hj��BR��B��H���Q�6�x   x   �!����������^��O���g8��P����^����������!��Ccg�xF��;'����c澈O��Ǡ��婏�0郾���/郾⩏�ʠ���O���c澔��;'�xF�=cg�x   x   ���k����Mſ@�Ͽ�$տ�$տ@�Ͽ�Mſi������ݪ��W7{�lT�0�/����<�u���V��穏�\��[��⩏�Q��q����<�
��3�/�oT�\7{�٪��x   x   �xʿ}�ݿ���2���u���2����~�ݿ�xʿd\���؜��L����]�g95�9����u���Ϡ��,w��eΌ�*w��ʠ��q������9�l95���]��L���؜�d\��x   x    ����r�
�Ȃ�ǂ�p�
������ڿ2���Ӥ�'-����b�M7�9��<꾃O��lj��=:��<:��hj���O���<�9�N7���b�(-���Ӥ�2����ڿx   x   &��sw�o��!�o��uw�'��x��5}�e�ǿt����؋���b�h95����c�?R��$����<��&���BR���c�
��l95���b��؋�t���`�ǿ6}�|��x   x   �:#��,��_1��_1��,��:#�&g�k����Eʿv���$-����]�1�/���H��yr��iޭ�gޭ�}r��B�ྔ�3�/���]�(-��t����Eʿ��j�&g�x   x   k6�[X>�aA�ZX>�k6� *�͈������`�ǿ�Ӥ��L��tT��;'�F����پ1I��uX��3I����پH���;'�oT��L���Ӥ�`�ǿ�����̈� *�x   x   W�F���L���L�U�F�n�;�},�͈�j�2}�2���؜�\7{�xF��Q�w���Ҿs��s���Ҿw���Q�xF�\7{��؜�2��6}�j�̈�},�m�;�x   x   g�R���U�h�R��I�m�;�*�&g�z����ڿf\��ߪ��Hcg�6�������(V̾={¾-V̾�����6�=cg�٪��d\����ڿ|��&g� *�m�;��I�x   